----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 25.12.2018 17:39:59
-- Design Name: 
-- Module Name: Snare - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_1164.ALL;


-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Snare is
    Port ( CLK : in STD_LOGIC;
           CE : in STD_LOGIC;
           RST : in STD_LOGIC;
           PLAY : in STD_LOGIC;
           SNARE_SAMP_O : out signed(7 downto 0)
           );
end Snare;

architecture Behavioral of Snare is

type memory is array (0 to 5551) of signed(7 downto 0);
constant snare_sound: memory := (
	x"08", x"12", x"14", x"1A", x"24", x"2E", x"2F", x"2F", x"2E", x"2B", x"25", x"28",
	x"26", x"1A", x"0E", x"07", x"FD", x"F9", x"FC", x"F6", x"FA", x"FD", x"FF", x"FD",
	x"FC", x"F1", x"E7", x"E3", x"DF", x"E1", x"DF", x"E0", x"DA", x"D7", x"D7", x"DD",
	x"E8", x"F5", x"FC", x"03", x"0D", x"0E", x"07", x"00", x"05", x"FF", x"0C", x"19",
	x"19", x"25", x"1C", x"27", x"22", x"0F", x"13", x"18", x"1E", x"1F", x"24", x"15",
	x"FF", x"F6", x"EE", x"F0", x"FA", x"FF", x"F9", x"F9", x"F6", x"EB", x"E5", x"EC",
	x"E5", x"E8", x"E7", x"E2", x"D1", x"C8", x"D6", x"CE", x"CF", x"D3", x"D4", x"DA",
	x"DB", x"E7", x"E2", x"E4", x"F3", x"FD", x"FF", x"0A", x"20", x"2D", x"35", x"3B",
	x"3E", x"36", x"43", x"52", x"46", x"4A", x"4B", x"4A", x"3E", x"3B", x"35", x"28",
	x"20", x"17", x"08", x"FC", x"EA", x"D0", x"C1", x"C0", x"C9", x"CD", x"CA", x"C2",
	x"C7", x"C3", x"BB", x"BE", x"C5", x"D0", x"D0", x"DB", x"CA", x"D0", x"D6", x"D8",
	x"EE", x"F7", x"F7", x"FD", x"24", x"17", x"24", x"3A", x"25", x"2C", x"27", x"2A",
	x"35", x"34", x"34", x"36", x"2C", x"32", x"31", x"2B", x"29", x"1D", x"24", x"16",
	x"08", x"FF", x"F4", x"ED", x"F0", x"F2", x"EB", x"F3", x"EE", x"E0", x"D5", x"C5",
	x"D7", x"D5", x"CD", x"BE", x"BF", x"CC", x"D9", x"F4", x"EF", x"EC", x"E5", x"EE",
	x"FD", x"0E", x"1D", x"0F", x"09", x"10", x"26", x"2E", x"1B", x"14", x"11", x"1C",
	x"21", x"17", x"0F", x"14", x"0F", x"16", x"21", x"21", x"16", x"0B", x"FF", x"0B",
	x"0B", x"10", x"17", x"FF", x"F7", x"F4", x"F0", x"E8", x"F3", x"E9", x"DC", x"DC",
	x"D5", x"C8", x"C3", x"C9", x"C6", x"D0", x"DA", x"F3", x"EB", x"E3", x"03", x"FD",
	x"13", x"24", x"1A", x"14", x"24", x"3D", x"24", x"2B", x"22", x"17", x"1A", x"15",
	x"F7", x"F4", x"05", x"FC", x"FC", x"0A", x"FD", x"ED", x"FC", x"00", x"FF", x"08",
	x"02", x"FB", x"F7", x"04", x"13", x"00", x"0C", x"00", x"EB", x"FD", x"FD", x"F9",
	x"00", x"E9", x"ED", x"F2", x"FB", x"F9", x"E0", x"E5", x"F1", x"05", x"09", x"08",
	x"ED", x"F0", x"01", x"0A", x"09", x"0E", x"17", x"0E", x"11", x"11", x"09", x"FE",
	x"0E", x"FB", x"05", x"13", x"14", x"0E", x"0C", x"06", x"F2", x"FF", x"FE", x"FE",
	x"F8", x"F5", x"EF", x"E8", x"F1", x"F5", x"E9", x"DF", x"E9", x"EF", x"F3", x"08",
	x"FC", x"F3", x"FB", x"F8", x"0C", x"03", x"10", x"0A", x"09", x"18", x"09", x"12",
	x"08", x"16", x"1D", x"13", x"11", x"09", x"0A", x"F5", x"FA", x"F9", x"EB", x"EC",
	x"DC", x"DB", x"EA", x"E2", x"E8", x"EC", x"EE", x"F0", x"F6", x"03", x"FC", x"02",
	x"04", x"0C", x"07", x"0E", x"00", x"F5", x"08", x"0D", x"0C", x"0C", x"12", x"09",
	x"01", x"03", x"10", x"10", x"10", x"0B", x"04", x"08", x"14", x"0F", x"F8", x"FE",
	x"FC", x"04", x"F9", x"07", x"FE", x"F4", x"FB", x"F6", x"FC", x"E9", x"F4", x"FB",
	x"EE", x"F8", x"04", x"FB", x"F4", x"ED", x"ED", x"F8", x"FC", x"F4", x"FC", x"F6",
	x"F0", x"F3", x"F7", x"FD", x"FF", x"08", x"08", x"04", x"10", x"11", x"0E", x"0A",
	x"0B", x"0D", x"0C", x"10", x"0E", x"10", x"15", x"19", x"0C", x"08", x"FD", x"F7",
	x"F5", x"F1", x"F7", x"F7", x"F4", x"EE", x"FB", x"F4", x"FB", x"F8", x"F2", x"FB",
	x"FA", x"F7", x"F3", x"F2", x"F2", x"F8", x"FC", x"FD", x"F0", x"FB", x"FA", x"F8",
	x"FF", x"F9", x"FB", x"F2", x"F5", x"FC", x"0A", x"09", x"11", x"0E", x"0D", x"0D",
	x"13", x"14", x"0C", x"11", x"0C", x"0B", x"0A", x"10", x"00", x"FB", x"FE", x"FC",
	x"08", x"06", x"FB", x"02", x"F7", x"FE", x"04", x"FA", x"F4", x"F5", x"F4", x"ED",
	x"F4", x"04", x"F3", x"F1", x"FA", x"FD", x"FB", x"FD", x"04", x"F0", x"F7", x"FD",
	x"F0", x"F2", x"FD", x"05", x"00", x"07", x"05", x"01", x"0B", x"0A", x"10", x"10",
	x"0E", x"10", x"04", x"FD", x"00", x"08", x"05", x"07", x"06", x"03", x"01", x"F9",
	x"FD", x"F7", x"F8", x"FF", x"FD", x"04", x"FE", x"FB", x"F4", x"F9", x"FC", x"00",
	x"FE", x"FA", x"FC", x"F7", x"F7", x"F7", x"F3", x"F2", x"EE", x"F4", x"01", x"F9",
	x"FA", x"01", x"FC", x"F9", x"FF", x"03", x"02", x"03", x"03", x"05", x"0A", x"0B",
	x"10", x"08", x"05", x"13", x"10", x"09", x"03", x"02", x"FC", x"FE", x"03", x"02",
	x"01", x"01", x"FB", x"01", x"FD", x"FB", x"FA", x"F8", x"08", x"FD", x"FA", x"FA",
	x"F5", x"F7", x"F8", x"FA", x"FA", x"FC", x"FD", x"FD", x"FE", x"F4", x"F8", x"F5",
	x"F8", x"02", x"00", x"00", x"FF", x"01", x"03", x"09", x"07", x"05", x"06", x"04",
	x"02", x"05", x"02", x"FF", x"05", x"FB", x"FD", x"05", x"03", x"0B", x"06", x"06",
	x"00", x"05", x"02", x"07", x"07", x"FC", x"FF", x"FD", x"01", x"F6", x"ED", x"EB",
	x"F4", x"F1", x"F2", x"FB", x"F6", x"FC", x"F7", x"F8", x"FE", x"FB", x"01", x"FE",
	x"03", x"02", x"04", x"09", x"02", x"07", x"05", x"04", x"02", x"01", x"06", x"01",
	x"04", x"FA", x"FB", x"FF", x"FD", x"04", x"FF", x"FE", x"03", x"FF", x"00", x"03",
	x"05", x"06", x"03", x"07", x"FF", x"06", x"00", x"FD", x"FA", x"F6", x"FA", x"F9",
	x"FF", x"F4", x"F0", x"F7", x"FC", x"01", x"FF", x"00", x"FC", x"FC", x"01", x"04",
	x"FD", x"02", x"05", x"FE", x"05", x"00", x"FD", x"FF", x"FA", x"FC", x"FE", x"02",
	x"FF", x"02", x"02", x"0A", x"0A", x"02", x"05", x"05", x"FF", x"04", x"06", x"03",
	x"00", x"00", x"05", x"FE", x"04", x"03", x"FB", x"FB", x"FB", x"FA", x"F9", x"FA",
	x"F4", x"F4", x"FA", x"F6", x"F8", x"F1", x"F6", x"F9", x"FE", x"02", x"FD", x"04",
	x"01", x"06", x"08", x"01", x"05", x"02", x"01", x"00", x"02", x"03", x"00", x"FD",
	x"01", x"FF", x"04", x"06", x"00", x"FD", x"FD", x"FE", x"FA", x"03", x"00", x"01",
	x"06", x"04", x"00", x"00", x"FD", x"FD", x"F7", x"FC", x"FF", x"FD", x"FF", x"FA",
	x"FC", x"FC", x"FF", x"00", x"08", x"07", x"07", x"00", x"00", x"05", x"FE", x"FF",
	x"00", x"FB", x"FE", x"FD", x"FB", x"FF", x"FB", x"00", x"FA", x"FE", x"00", x"00",
	x"FE", x"00", x"FD", x"FB", x"FB", x"FD", x"06", x"03", x"03", x"02", x"04", x"06",
	x"07", x"04", x"FF", x"FF", x"00", x"01", x"FC", x"FB", x"F7", x"FA", x"FA", x"00",
	x"02", x"FE", x"00", x"FC", x"FF", x"FA", x"02", x"FD", x"FB", x"FC", x"F9", x"00",
	x"FF", x"FE", x"F9", x"FB", x"01", x"FF", x"03", x"00", x"00", x"01", x"04", x"00",
	x"00", x"04", x"04", x"07", x"08", x"06", x"FF", x"03", x"FF", x"FA", x"04", x"FE",
	x"FE", x"F9", x"FF", x"01", x"F8", x"FE", x"FB", x"FB", x"01", x"FE", x"FE", x"FC",
	x"FC", x"FB", x"F9", x"FC", x"FE", x"01", x"02", x"05", x"01", x"FE", x"05", x"03",
	x"03", x"03", x"01", x"FF", x"FC", x"FA", x"F9", x"F7", x"FE", x"03", x"00", x"05",
	x"02", x"03", x"02", x"00", x"FE", x"FB", x"01", x"FD", x"FD", x"FF", x"F9", x"FC",
	x"F9", x"F9", x"FD", x"FE", x"02", x"02", x"03", x"FE", x"FE", x"02", x"00", x"04",
	x"02", x"08", x"02", x"04", x"01", x"FE", x"FF", x"FF", x"FE", x"FF", x"03", x"FC",
	x"FE", x"FB", x"F9", x"FB", x"FC", x"01", x"FC", x"FD", x"FC", x"F9", x"FD", x"FF",
	x"FB", x"02", x"03", x"00", x"03", x"01", x"00", x"02", x"01", x"03", x"02", x"03",
	x"FF", x"FC", x"F9", x"FC", x"FB", x"01", x"FF", x"01", x"04", x"02", x"03", x"04",
	x"00", x"FD", x"FF", x"FE", x"02", x"00", x"FC", x"F9", x"F9", x"F9", x"F9", x"F6",
	x"FD", x"01", x"07", x"05", x"FF", x"FD", x"FE", x"03", x"03", x"03", x"04", x"05",
	x"02", x"FE", x"01", x"00", x"FF", x"00", x"03", x"FF", x"01", x"00", x"FA", x"FB",
	x"FC", x"FB", x"FC", x"FE", x"FF", x"FE", x"01", x"FE", x"FE", x"FF", x"00", x"FF",
	x"FE", x"FE", x"01", x"FF", x"03", x"FB", x"FB", x"FF", x"FF", x"00", x"02", x"04",
	x"FF", x"01", x"FD", x"FD", x"FE", x"FF", x"01", x"01", x"03", x"00", x"00", x"FF",
	x"FD", x"02", x"FE", x"FE", x"00", x"F7", x"FB", x"F6", x"F8", x"FE", x"00", x"FE",
	x"01", x"02", x"02", x"05", x"03", x"03", x"06", x"05", x"01", x"FD", x"FE", x"00",
	x"FD", x"00", x"FC", x"00", x"00", x"03", x"03", x"00", x"FD", x"FC", x"FC", x"FD",
	x"FD", x"FD", x"FC", x"FF", x"FF", x"02", x"FF", x"FD", x"FE", x"FF", x"03", x"03",
	x"03", x"01", x"FA", x"FE", x"FD", x"FD", x"FF", x"01", x"00", x"00", x"FF", x"00",
	x"01", x"01", x"01", x"FC", x"FF", x"00", x"FF", x"FE", x"FF", x"FD", x"FC", x"00",
	x"00", x"FD", x"FD", x"FC", x"FA", x"FC", x"FD", x"FF", x"FD", x"FE", x"00", x"01",
	x"04", x"04", x"05", x"03", x"02", x"05", x"03", x"01", x"02", x"00", x"FD", x"FC",
	x"FC", x"FD", x"FE", x"FC", x"01", x"FE", x"01", x"FE", x"FE", x"FE", x"FA", x"FD",
	x"FC", x"F9", x"00", x"01", x"FC", x"FF", x"FF", x"01", x"01", x"FF", x"02", x"FE",
	x"00", x"FF", x"FC", x"FE", x"02", x"01", x"00", x"00", x"01", x"01", x"00", x"FF",
	x"01", x"FD", x"01", x"00", x"FF", x"FF", x"FA", x"FE", x"FD", x"FE", x"FD", x"FF",
	x"FF", x"FE", x"FF", x"FD", x"FC", x"FD", x"FF", x"00", x"00", x"FE", x"FF", x"01",
	x"02", x"02", x"02", x"06", x"03", x"01", x"FF", x"FC", x"F9", x"FD", x"FD", x"FE",
	x"FE", x"00", x"00", x"FF", x"FE", x"FE", x"FC", x"00", x"01", x"FD", x"01", x"FF",
	x"FF", x"FC", x"FC", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"02", x"00",
	x"FF", x"01", x"00", x"01", x"00", x"01", x"FD", x"FD", x"FB", x"FF", x"00", x"01",
	x"04", x"01", x"FF", x"FD", x"FD", x"FA", x"FA", x"FB", x"FD", x"FE", x"FE", x"00",
	x"FF", x"FE", x"01", x"00", x"01", x"01", x"01", x"00", x"02", x"01", x"01", x"01",
	x"04", x"03", x"02", x"01", x"02", x"FD", x"FD", x"FE", x"FB", x"FA", x"00", x"FD",
	x"FD", x"01", x"FE", x"FB", x"FE", x"00", x"FF", x"04", x"02", x"00", x"FF", x"FC",
	x"FD", x"FA", x"FE", x"FD", x"FE", x"01", x"01", x"00", x"02", x"01", x"00", x"01",
	x"02", x"00", x"00", x"FD", x"FE", x"FD", x"FD", x"FF", x"02", x"00", x"03", x"01",
	x"FE", x"FF", x"FC", x"FC", x"FB", x"FC", x"FC", x"FE", x"FF", x"01", x"FC", x"FF",
	x"00", x"01", x"02", x"03", x"00", x"04", x"03", x"01", x"02", x"FE", x"FE", x"FE",
	x"FF", x"03", x"00", x"00", x"FF", x"FF", x"FC", x"FD", x"FD", x"FB", x"FF", x"FD",
	x"FE", x"FD", x"FE", x"01", x"00", x"00", x"01", x"02", x"00", x"FD", x"FC", x"F9",
	x"FD", x"FE", x"00", x"01", x"01", x"FF", x"02", x"03", x"00", x"02", x"01", x"00",
	x"02", x"00", x"FE", x"FF", x"FB", x"FE", x"FF", x"FD", x"00", x"00", x"FE", x"00",
	x"00", x"FE", x"FE", x"FD", x"FE", x"FE", x"FC", x"FF", x"FE", x"FE", x"FE", x"FF",
	x"FE", x"03", x"03", x"02", x"02", x"00", x"FD", x"FC", x"FD", x"00", x"FD", x"02",
	x"02", x"02", x"FF", x"FF", x"FD", x"FD", x"FD", x"00", x"FF", x"FD", x"FD", x"FD",
	x"01", x"01", x"02", x"01", x"FF", x"FE", x"00", x"FF", x"FE", x"FB", x"FE", x"FE",
	x"FF", x"00", x"02", x"FD", x"FD", x"00", x"FE", x"01", x"04", x"03", x"01", x"00",
	x"FE", x"FD", x"FB", x"FA", x"FC", x"FC", x"FE", x"00", x"FF", x"FF", x"FE", x"FD",
	x"01", x"01", x"01", x"01", x"FD", x"FD", x"FD", x"FD", x"FF", x"01", x"01", x"01",
	x"04", x"04", x"03", x"00", x"FD", x"FF", x"FD", x"FE", x"FF", x"00", x"01", x"FF",
	x"FC", x"FE", x"00", x"FF", x"FF", x"01", x"FF", x"02", x"01", x"FF", x"FC", x"FE",
	x"FE", x"FF", x"00", x"FD", x"FE", x"FC", x"FD", x"FD", x"FF", x"FE", x"FF", x"FF",
	x"00", x"FE", x"FD", x"FD", x"FE", x"01", x"02", x"04", x"05", x"03", x"00", x"FF",
	x"FE", x"FB", x"FD", x"FF", x"FC", x"FC", x"00", x"FE", x"FE", x"00", x"03", x"FF",
	x"02", x"00", x"FE", x"FF", x"FD", x"FB", x"FF", x"FE", x"FF", x"01", x"01", x"00",
	x"01", x"00", x"01", x"01", x"00", x"00", x"02", x"FD", x"FD", x"FD", x"FC", x"FE",
	x"FF", x"FE", x"00", x"03", x"03", x"02", x"00", x"00", x"FE", x"FC", x"FC", x"FD",
	x"FD", x"FF", x"FD", x"FE", x"FD", x"00", x"FF", x"01", x"FE", x"01", x"00", x"FF",
	x"01", x"FE", x"FF", x"04", x"03", x"02", x"02", x"00", x"00", x"FE", x"FD", x"FD",
	x"FF", x"00", x"FF", x"00", x"FE", x"FD", x"FD", x"FE", x"FE", x"02", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FC", x"FD", x"FF", x"FF", x"FE", x"FF", x"FD", x"FF",
	x"00", x"00", x"01", x"03", x"00", x"FF", x"FE", x"FA", x"FD", x"FE", x"FE", x"FE",
	x"FF", x"03", x"04", x"02", x"02", x"FD", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE",
	x"00", x"FE", x"FF", x"00", x"00", x"FF", x"02", x"01", x"02", x"01", x"00", x"FF",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FD", x"FE", x"FD", x"FE", x"FF", x"00",
	x"01", x"FE", x"FD", x"FD", x"FE", x"FC", x"FE", x"01", x"01", x"00", x"01", x"00",
	x"FF", x"FF", x"00", x"FB", x"FD", x"FF", x"FE", x"00", x"00", x"FF", x"00", x"01",
	x"02", x"02", x"03", x"00", x"FF", x"FC", x"FD", x"FF", x"FD", x"FE", x"FF", x"01",
	x"FF", x"FF", x"00", x"FE", x"FF", x"FE", x"00", x"00", x"FF", x"FC", x"FF", x"FB",
	x"FC", x"FC", x"FD", x"FF", x"01", x"02", x"03", x"01", x"02", x"FF", x"01", x"FF",
	x"FE", x"FE", x"FD", x"FE", x"FF", x"FE", x"FE", x"00", x"FF", x"04", x"03", x"01",
	x"FF", x"FD", x"FF", x"FD", x"FC", x"FF", x"00", x"01", x"02", x"FE", x"FF", x"FF",
	x"FE", x"00", x"FD", x"FF", x"FD", x"00", x"FF", x"FC", x"FC", x"01", x"03", x"01",
	x"02", x"01", x"FF", x"00", x"FF", x"FE", x"FF", x"FE", x"FC", x"FE", x"FE", x"FD",
	x"FD", x"FE", x"00", x"FE", x"02", x"01", x"01", x"FE", x"FE", x"FA", x"FD", x"FE",
	x"FE", x"01", x"01", x"01", x"02", x"02", x"03", x"00", x"FE", x"FF", x"FF", x"00",
	x"00", x"FC", x"FC", x"FD", x"FD", x"FF", x"01", x"01", x"01", x"FF", x"FF", x"00",
	x"FE", x"00", x"00", x"FF", x"FF", x"01", x"FD", x"FE", x"FF", x"FD", x"FF", x"FF",
	x"00", x"00", x"01", x"FE", x"FF", x"FE", x"FE", x"FE", x"00", x"00", x"FF", x"02",
	x"02", x"00", x"01", x"FF", x"FE", x"FE", x"FE", x"FF", x"FE", x"FB", x"FE", x"FD",
	x"FE", x"FF", x"01", x"03", x"FF", x"FF", x"FF", x"FC", x"FE", x"FD", x"FE", x"FF",
	x"01", x"FF", x"02", x"02", x"FF", x"00", x"FF", x"01", x"00", x"01", x"00", x"FD",
	x"FF", x"FD", x"FD", x"FD", x"FD", x"FF", x"01", x"01", x"00", x"01", x"FF", x"00",
	x"00", x"00", x"00", x"FD", x"FE", x"FC", x"FB", x"FD", x"FD", x"00", x"01", x"03",
	x"02", x"00", x"FF", x"FF", x"FF", x"FD", x"00", x"00", x"00", x"02", x"FF", x"00",
	x"00", x"00", x"FF", x"00", x"FE", x"00", x"FE", x"FD", x"FC", x"FF", x"FE", x"FF",
	x"00", x"FE", x"FE", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"01", x"FF",
	x"FF", x"FD", x"FE", x"FF", x"00", x"FF", x"01", x"FF", x"01", x"00", x"FE", x"FD",
	x"FB", x"FE", x"FC", x"FF", x"02", x"FF", x"01", x"00", x"00", x"00", x"FF", x"00",
	x"FE", x"FF", x"FD", x"FD", x"FF", x"FC", x"FF", x"FF", x"01", x"01", x"02", x"02",
	x"02", x"00", x"00", x"01", x"01", x"FF", x"01", x"FF", x"00", x"FF", x"FB", x"FE",
	x"FE", x"00", x"FD", x"FF", x"FD", x"FF", x"00", x"FE", x"FE", x"FD", x"FC", x"FF",
	x"FF", x"01", x"00", x"FF", x"01", x"01", x"01", x"FE", x"00", x"FD", x"FD", x"FD",
	x"FF", x"FF", x"FF", x"01", x"FF", x"00", x"02", x"02", x"00", x"FF", x"FE", x"FD",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"01", x"00", x"FE", x"FE", x"FF",
	x"FF", x"FD", x"FD", x"FC", x"FD", x"00", x"FF", x"00", x"01", x"00", x"01", x"01",
	x"03", x"03", x"01", x"01", x"01", x"FF", x"FC", x"FC", x"FB", x"FD", x"FF", x"FE",
	x"FF", x"00", x"00", x"01", x"00", x"FF", x"FD", x"FD", x"FF", x"00", x"FF", x"FF",
	x"FF", x"00", x"01", x"00", x"00", x"00", x"01", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FE", x"00", x"FF", x"01", x"00", x"FD", x"FE", x"FD", x"00", x"FE", x"FF",
	x"FF", x"FE", x"00", x"FE", x"FF", x"FE", x"00", x"00", x"FF", x"01", x"00", x"FF",
	x"00", x"FE", x"FE", x"FD", x"FE", x"FE", x"00", x"01", x"02", x"00", x"04", x"02",
	x"02", x"01", x"00", x"FF", x"FD", x"FC", x"FD", x"FC", x"FE", x"FE", x"FF", x"FF",
	x"00", x"00", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"FF", x"FF", x"FE", x"FD",
	x"FF", x"FF", x"FE", x"00", x"00", x"01", x"00", x"01", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FD", x"00", x"01", x"00", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FD", x"FC", x"FE", x"FF", x"00", x"01", x"00", x"00", x"FE", x"FF",
	x"FF", x"FD", x"FE", x"FF", x"FE", x"00", x"00", x"01", x"01", x"00", x"02", x"FF",
	x"00", x"FD", x"FE", x"FD", x"FE", x"FD", x"FD", x"FD", x"FF", x"01", x"00", x"01",
	x"FF", x"01", x"01", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FD", x"FE", x"FC",
	x"FD", x"00", x"01", x"01", x"02", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FE",
	x"FD", x"FF", x"FE", x"00", x"FF", x"FF", x"FF", x"01", x"FF", x"00", x"FF", x"FD",
	x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"00", x"FE", x"00", x"00", x"01", x"FF",
	x"FF", x"02", x"00", x"00", x"FF", x"FE", x"FF", x"00", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FD", x"FF", x"FE", x"FD", x"FF", x"FF", x"FD", x"00", x"01", x"00",
	x"00", x"01", x"02", x"02", x"02", x"FF", x"FC", x"FC", x"FB", x"FD", x"FD", x"FF",
	x"00", x"00", x"01", x"00", x"FF", x"FF", x"01", x"01", x"01", x"00", x"FE", x"00",
	x"FE", x"FD", x"FE", x"FE", x"00", x"01", x"00", x"00", x"FE", x"FE", x"FF", x"00",
	x"FE", x"FF", x"FC", x"FD", x"FD", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"01",
	x"02", x"01", x"00", x"FF", x"FF", x"FD", x"FE", x"FD", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FE", x"FF", x"FE", x"FF", x"00", x"FE", x"00", x"00", x"FF",
	x"FF", x"01", x"01", x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"00", x"FE", x"FF",
	x"FF", x"00", x"FF", x"01", x"01", x"02", x"01", x"01", x"FF", x"00", x"FE", x"FE",
	x"FE", x"FE", x"FD", x"FF", x"FF", x"01", x"00", x"00", x"FF", x"00", x"00", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FF", x"FF", x"FE", x"01", x"00", x"01", x"00", x"00",
	x"00", x"FF", x"FD", x"FE", x"FC", x"FE", x"FF", x"FF", x"00", x"FE", x"00", x"FE",
	x"FF", x"01", x"FF", x"00", x"01", x"FF", x"00", x"FD", x"00", x"FF", x"FE", x"01",
	x"FE", x"FE", x"FE", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"00", x"01", x"01", x"01", x"03", x"00", x"FF", x"FE", x"FC", x"FD", x"FD",
	x"FD", x"FE", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"01", x"FE",
	x"FF", x"FF", x"FE", x"00", x"FE", x"FF", x"00", x"01", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FE", x"FF", x"FD", x"FF", x"FF", x"01",
	x"00", x"01", x"00", x"00", x"FF", x"FF", x"FC", x"FD", x"FE", x"FE", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"01", x"01", x"01", x"FF", x"01", x"00", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF",
	x"FD", x"FE", x"FD", x"00", x"FE", x"00", x"01", x"00", x"01", x"00", x"00", x"FD",
	x"FF", x"FC", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"01", x"00", x"01",
	x"02", x"01", x"FF", x"FF", x"FD", x"FD", x"FD", x"FE", x"FE", x"FC", x"FE", x"FE",
	x"00", x"FF", x"FF", x"00", x"00", x"01", x"FF", x"00", x"FF", x"FF", x"00", x"FF",
	x"01", x"FF", x"FE", x"FF", x"FF", x"FE", x"00", x"FE", x"00", x"FE", x"FF", x"FE",
	x"FD", x"FE", x"FF", x"00", x"00", x"02", x"00", x"01", x"01", x"FF", x"00", x"FE",
	x"FF", x"FF", x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"FF", x"01", x"FF",
	x"00", x"00", x"FE", x"FF", x"FE", x"FE", x"FD", x"FF", x"FF", x"00", x"01", x"FF",
	x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"01", x"02", x"02", x"00", x"01", x"FF", x"FF", x"00", x"FD", x"FF", x"FF",
	x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FD", x"FE", x"FF", x"01", x"00", x"01", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"FF", x"01",
	x"00", x"FF", x"FF", x"FD", x"FF", x"FD", x"00", x"FE", x"FF", x"FE", x"00", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"00", x"01", x"02", x"01", x"01", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"00", x"00", x"00", x"00", x"01", x"00", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"00", x"FE", x"00", x"FF",
	x"FE", x"FE", x"FD", x"FF", x"FE", x"00", x"FF", x"01", x"01", x"00", x"01", x"00",
	x"FF", x"FE", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FF", x"00", x"00", x"00",
	x"00", x"01", x"00", x"01", x"FE", x"FF", x"FE", x"FE", x"00", x"FF", x"01", x"00",
	x"01", x"00", x"01", x"FE", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FC", x"FE",
	x"FD", x"FE", x"FF", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"01", x"FF",
	x"FF", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"00", x"FF", x"01", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"00", x"FE", x"FF", x"FD", x"FD", x"FF", x"FF", x"00", x"FF", x"01",
	x"FF", x"FF", x"00", x"FE", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FE",
	x"FF", x"FF", x"01", x"FF", x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FC", x"FE",
	x"FF", x"FF", x"01", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FD",
	x"FE", x"FD", x"FE", x"FE", x"FE", x"00", x"FF", x"01", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FD", x"FF", x"FF", x"00", x"FF",
	x"00", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"01",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"00", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"01", x"FF", x"00", x"00", x"FE", x"FE", x"FD", x"FF", x"FE", x"00",
	x"00", x"00", x"01", x"01", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FE", x"FE",
	x"FE", x"FD", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"00", x"01", x"FF", x"00",
	x"FF", x"00", x"FE", x"FE", x"FE", x"FC", x"FE", x"FE", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FE", x"01", x"FF", x"00", x"FE", x"FF", x"FD", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"01", x"FF", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FE", x"00", x"FE", x"00", x"00", x"FF", x"00", x"FE", x"FE", x"FD", x"FD",
	x"FE", x"FE", x"FF", x"00", x"00", x"FF", x"01", x"00", x"01", x"01", x"01", x"00",
	x"FF", x"FF", x"FC", x"FE", x"FD", x"FE", x"FF", x"00", x"00", x"01", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FD", x"FE", x"FC", x"FE", x"FF", x"00", x"FF",
	x"00", x"00", x"FE", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FD", x"FF", x"FE", x"01", x"00", x"00", x"FE", x"FF", x"FD", x"FF", x"FF", x"FD",
	x"FF", x"FE", x"01", x"FF", x"00", x"00", x"00", x"01", x"FF", x"00", x"00", x"FE",
	x"FF", x"FF", x"FD", x"FE", x"FE", x"00", x"FF", x"FE", x"00", x"FF", x"01", x"00",
	x"FF", x"01", x"FF", x"FF", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FE",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"02", x"00", x"00",
	x"FF", x"00", x"FE", x"FF", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF",
	x"00", x"FF", x"01", x"FF", x"FF", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"00",
	x"FF", x"01", x"FE", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FE", x"00", x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FE", x"FF", x"FD", x"FE", x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"00",
	x"00", x"01", x"00", x"00", x"00", x"00", x"FE", x"FF", x"FD", x"FF", x"FE", x"FF",
	x"FE", x"00", x"FF", x"00", x"00", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FD", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"00", x"FF", x"01", x"FF", x"00",
	x"00", x"FE", x"FE", x"FD", x"FF", x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"02",
	x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"00", x"00", x"FF", x"01", x"FF", x"00", x"00", x"FE", x"00", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"01", x"00", x"00",
	x"FE", x"00", x"FE", x"FF", x"FF", x"FE", x"00", x"FE", x"00", x"FF", x"00", x"FE",
	x"00", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"01", x"01", x"FF",
	x"00", x"FF", x"00", x"FE", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE",
	x"FF", x"FE", x"FD", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"01", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FE", x"FF",
	x"FF", x"00", x"01", x"00", x"01", x"FF", x"00", x"00", x"FF", x"FE", x"FE", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FD", x"FF", x"FE", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"00", x"FE", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FE", x"00", x"00",
	x"01", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"00", x"FE", x"00", x"00", x"FF", x"00", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FE", x"FE", x"FD", x"FE", x"FD", x"FF", x"FF", x"FF", x"01", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"00", x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"00", x"FE", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FE", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"00", x"FF", x"FF", x"FE", x"FF", x"00", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"00", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"00", x"FE", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FE", x"00", x"01",
	x"00", x"01", x"01", x"01", x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"00",
	x"00", x"FE", x"00", x"FF", x"FF", x"FE", x"00", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF",
	x"01", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FD", x"FF",
	x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FE", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FE", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FE", x"00",
	x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"00", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FE", x"00",
	x"FF", x"00", x"FF", x"00", x"FE", x"00", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF",
	x"FE", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FE", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FE", x"00", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FE", x"00", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"FE", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"00", x"00", x"00", x"00",
	x"FE", x"00", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00",
	x"FE", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"FE", x"FF", x"FE",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"00", x"FE", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"FE", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FE", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"00",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"00", x"FF", x"FE", x"00", x"FE", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"00",
	x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"00",
	x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"00", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"FF", x"FE", x"00", x"FF",
	x"00", x"FF", x"FF", x"FE", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FE", x"00",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"00",
	x"FF", x"00", x"FE", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FE", x"00", x"FE", x"00", x"FF", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"FE", x"00", x"FE", x"FF", x"FF", x"00", x"FE",
	x"FF", x"00", x"FF", x"FF", x"00", x"FE", x"FE", x"FF", x"FE", x"FF", x"FE", x"00",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"00", x"FF", x"00", x"00", x"FE", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"00", x"FF", x"FF", x"FF", x"FE",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FE", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FE", x"00", x"FE", x"FF", x"FE",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FE",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FE",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"FE", x"00", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF"
	);
	
signal cnt_out: integer := 0;	
signal play_sound: std_logic := '0';
constant cnt_max: integer := 5551;
signal out_signal: signed(7 downto 0) := x"00";

begin
	
process (CLK)
begin
    if rising_edge(CLK) then
        if RST = '1' then
            play_sound <= '0';
        elsif PLAY = '1' then
            play_sound <= '1';
        elsif PLAY = '0' and cnt_out = cnt_max then
            play_sound <= '0';
        end if;
    end if;
end process;

	
-- 12bit counter
process (CLK)
begin     
    if rising_edge(CLK) then
        if RST = '1' then
            cnt_out <= 0;
        elsif CE = '1' and play_sound = '1' then
            cnt_out <= cnt_out + 1;       
        end if;
        if cnt_out = cnt_max then
            cnt_out <= 0;            
        end if;        
    end if;
end process;

process (CLK) 
begin
    if rising_edge(CLK) then
        if RST = '1' then
            out_signal <= x"00";
        elsif CE = '1' then
            out_signal <= snare_sound(cnt_out);
        end if;
    end if;    
end process;

SNARE_SAMP_O <= out_signal;

end Behavioral;