----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 22.12.2018 23:25:25
-- Design Name: 
-- Module Name: Kick - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_1164.ALL;


-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Kick is
    Port ( CLK : in STD_LOGIC;
           CE : in STD_LOGIC;
           RST : in STD_LOGIC;
           PLAY : in STD_LOGIC;
           KICK_SAMP_O : out signed(7 downto 0)
           );
end Kick;

architecture Behavioral of Kick is

type memory is array (0 to 9557) of signed(7 downto 0);
constant kick_sound: memory := (
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"02", x"04", x"05", x"06", x"06", x"07", x"07", x"07", x"08", x"08", x"09", x"09",
	x"08", x"08", x"07", x"07", x"08", x"0A", x"0C", x"0F", x"11", x"12", x"13", x"14",
	x"16", x"16", x"17", x"17", x"17", x"16", x"16", x"15", x"15", x"16", x"18", x"19",
	x"19", x"1A", x"1B", x"1D", x"1F", x"22", x"23", x"23", x"22", x"22", x"22", x"21",
	x"20", x"1F", x"1F", x"1E", x"1D", x"1D", x"1D", x"1E", x"1F", x"21", x"22", x"23",
	x"24", x"24", x"24", x"23", x"21", x"20", x"22", x"22", x"1E", x"1C", x"1E", x"21",
	x"20", x"1E", x"1D", x"20", x"25", x"24", x"1F", x"1A", x"1D", x"25", x"2C", x"29",
	x"20", x"1B", x"1F", x"27", x"2B", x"28", x"21", x"1B", x"1A", x"1D", x"22", x"27",
	x"28", x"24", x"1D", x"17", x"15", x"19", x"22", x"2A", x"2D", x"27", x"19", x"10",
	x"0F", x"17", x"21", x"28", x"29", x"23", x"17", x"0E", x"0B", x"11", x"19", x"23",
	x"2C", x"2C", x"25", x"19", x"13", x"15", x"18", x"1B", x"1E", x"20", x"20", x"1F",
	x"1F", x"23", x"25", x"1F", x"13", x"06", x"03", x"0C", x"1A", x"27", x"30", x"36",
	x"37", x"31", x"29", x"23", x"1F", x"1C", x"18", x"12", x"0A", x"FF", x"F2", x"EA",
	x"ED", x"F6", x"03", x"0F", x"10", x"09", x"FB", x"E8", x"D5", x"C9", x"C2", x"C3",
	x"C7", x"CC", x"D1", x"D7", x"DC", x"E0", x"E4", x"E7", x"E8", x"EB", x"ED", x"F0",
	x"F1", x"F1", x"F1", x"EE", x"E8", x"DE", x"D5", x"D3", x"D6", x"DA", x"DB", x"D6",
	x"D0", x"CC", x"CA", x"CA", x"CD", x"CE", x"CF", x"D1", x"D0", x"CD", x"CE", x"D3",
	x"D1", x"C9", x"BD", x"B1", x"A7", x"9F", x"9B", x"99", x"99", x"9B", x"9E", x"A4",
	x"A9", x"AB", x"AD", x"B2", x"BB", x"BD", x"BD", x"B8", x"AE", x"A2", x"98", x"94",
	x"93", x"92", x"8D", x"88", x"85", x"84", x"86", x"8A", x"90", x"96", x"9D", x"A1",
	x"A0", x"9E", x"9C", x"9D", x"9E", x"A2", x"A8", x"B0", x"B6", x"BA", x"BA", x"B2",
	x"A6", x"9F", x"9C", x"9C", x"9B", x"99", x"96", x"94", x"98", x"9D", x"A3", x"A7",
	x"AB", x"B0", x"B4", x"B6", x"B5", x"B4", x"B3", x"B3", x"B3", x"B3", x"B5", x"B9",
	x"BA", x"B9", x"B9", x"B8", x"B7", x"B4", x"B0", x"AF", x"B0", x"AE", x"AA", x"A4",
	x"9D", x"96", x"95", x"9C", x"A1", x"A2", x"A5", x"A7", x"AB", x"B1", x"B8", x"C1",
	x"C9", x"D1", x"D7", x"DB", x"DC", x"DA", x"D5", x"CD", x"C8", x"C3", x"BE", x"BB",
	x"BC", x"BE", x"C0", x"C1", x"C4", x"C9", x"CF", x"D6", x"D8", x"DB", x"E1", x"EB",
	x"F4", x"F8", x"F7", x"F6", x"F4", x"F1", x"EF", x"F1", x"F4", x"F8", x"FE", x"04",
	x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"0A", x"10", x"1A", x"24", x"2C",
	x"30", x"30", x"2B", x"25", x"21", x"20", x"20", x"23", x"27", x"28", x"29", x"2C",
	x"31", x"38", x"3F", x"41", x"40", x"3E", x"3B", x"36", x"32", x"31", x"32", x"33",
	x"32", x"33", x"39", x"42", x"4C", x"56", x"5E", x"63", x"64", x"62", x"61", x"61",
	x"63", x"64", x"65", x"65", x"62", x"60", x"5F", x"61", x"63", x"66", x"66", x"65",
	x"64", x"64", x"62", x"62", x"65", x"6E", x"79", x"7E", x"7C", x"7C", x"7C", x"7C",
	x"7C", x"7C", x"7D", x"7D", x"7C", x"7B", x"7A", x"79", x"7A", x"7B", x"7A", x"7B",
	x"7A", x"7A", x"7B", x"7B", x"7A", x"77", x"74", x"71", x"6F", x"6C", x"69", x"67",
	x"68", x"6C", x"71", x"75", x"79", x"7B", x"7C", x"7C", x"77", x"6E", x"64", x"5E",
	x"5C", x"5F", x"64", x"69", x"6E", x"70", x"70", x"70", x"6F", x"6F", x"6F", x"70",
	x"70", x"6F", x"6E", x"6F", x"6F", x"6E", x"6A", x"66", x"64", x"63", x"62", x"61",
	x"5F", x"5E", x"5E", x"5F", x"60", x"5F", x"5E", x"5E", x"5E", x"5E", x"5B", x"58",
	x"57", x"59", x"5C", x"60", x"65", x"68", x"68", x"66", x"63", x"63", x"64", x"64",
	x"63", x"61", x"60", x"5E", x"5C", x"59", x"55", x"50", x"4E", x"49", x"43", x"40",
	x"40", x"43", x"47", x"49", x"47", x"45", x"44", x"45", x"45", x"46", x"45", x"44",
	x"42", x"3F", x"39", x"32", x"2B", x"28", x"28", x"2A", x"2B", x"2C", x"29", x"27",
	x"26", x"24", x"23", x"22", x"21", x"1C", x"15", x"0E", x"07", x"03", x"00", x"00",
	x"02", x"03", x"07", x"0D", x"13", x"15", x"12", x"0F", x"0E", x"0E", x"0F", x"0E",
	x"0C", x"0A", x"08", x"08", x"06", x"03", x"FF", x"FC", x"FC", x"FD", x"FD", x"FC",
	x"FA", x"F9", x"F6", x"F3", x"EF", x"EB", x"E6", x"E5", x"E6", x"E9", x"EC", x"EA",
	x"E8", x"E4", x"E2", x"E3", x"E5", x"E8", x"EA", x"EA", x"E8", x"E2", x"DD", x"D9",
	x"D8", x"D8", x"D6", x"D1", x"CC", x"CB", x"CA", x"C9", x"C6", x"C4", x"C3", x"C3",
	x"BF", x"B9", x"B1", x"AC", x"AA", x"AB", x"AD", x"B1", x"B3", x"B3", x"B1", x"B0",
	x"AD", x"AA", x"A7", x"A4", x"A5", x"A7", x"AA", x"AB", x"AB", x"AB", x"AB", x"AB",
	x"AB", x"AA", x"A8", x"A5", x"A2", x"9D", x"9B", x"9C", x"9F", x"A3", x"A5", x"A7",
	x"A8", x"A9", x"A7", x"A5", x"A3", x"A2", x"A3", x"A3", x"A1", x"9D", x"98", x"92",
	x"8C", x"86", x"83", x"85", x"88", x"8C", x"8E", x"8E", x"8E", x"8C", x"8C", x"8C",
	x"8C", x"89", x"87", x"86", x"87", x"89", x"8C", x"8E", x"90", x"93", x"95", x"96",
	x"95", x"94", x"94", x"96", x"97", x"96", x"91", x"8B", x"87", x"86", x"87", x"89",
	x"8B", x"8D", x"8E", x"8F", x"8E", x"8F", x"92", x"93", x"91", x"8E", x"8C", x"8A",
	x"89", x"88", x"88", x"8A", x"8D", x"91", x"96", x"97", x"98", x"98", x"97", x"95",
	x"91", x"8B", x"87", x"85", x"84", x"84", x"86", x"88", x"88", x"89", x"8B", x"8D",
	x"8E", x"8E", x"8F", x"8F", x"8E", x"8F", x"8F", x"90", x"93", x"94", x"94", x"94",
	x"93", x"92", x"92", x"92", x"93", x"95", x"95", x"92", x"8F", x"8D", x"8D", x"8E",
	x"8F", x"90", x"91", x"94", x"95", x"95", x"95", x"95", x"95", x"93", x"91", x"8D",
	x"89", x"87", x"88", x"8B", x"90", x"93", x"96", x"98", x"9B", x"9B", x"99", x"97",
	x"97", x"9A", x"9F", x"A4", x"A6", x"A6", x"A4", x"A0", x"9E", x"9F", x"A2", x"A5",
	x"A8", x"A8", x"A6", x"A5", x"A4", x"A5", x"A9", x"AC", x"AF", x"B1", x"B0", x"AF",
	x"AF", x"B0", x"B1", x"B2", x"B4", x"B6", x"B9", x"BC", x"BD", x"BF", x"BF", x"BE",
	x"BC", x"BB", x"BB", x"BD", x"C2", x"C8", x"CF", x"D5", x"D9", x"DB", x"DC", x"DC",
	x"DC", x"DC", x"DA", x"D7", x"D3", x"CF", x"CC", x"CB", x"C9", x"CB", x"D0", x"D6",
	x"DD", x"E4", x"E8", x"EB", x"ED", x"ED", x"EC", x"EB", x"EB", x"EC", x"EE", x"F1",
	x"F6", x"FC", x"01", x"02", x"01", x"01", x"04", x"0A", x"10", x"13", x"15", x"16",
	x"16", x"17", x"17", x"17", x"19", x"1E", x"25", x"2D", x"31", x"33", x"33", x"32",
	x"32", x"34", x"35", x"35", x"34", x"34", x"36", x"38", x"39", x"3B", x"3E", x"40",
	x"41", x"41", x"42", x"42", x"43", x"44", x"46", x"48", x"4A", x"4C", x"4C", x"4C",
	x"4B", x"49", x"47", x"44", x"44", x"44", x"44", x"46", x"4A", x"50", x"55", x"5A",
	x"5E", x"60", x"5E", x"5C", x"5B", x"59", x"5A", x"5C", x"5C", x"5D", x"5F", x"61",
	x"65", x"69", x"69", x"66", x"64", x"65", x"67", x"66", x"65", x"64", x"63", x"62",
	x"60", x"5D", x"5B", x"5B", x"5C", x"5E", x"62", x"68", x"6D", x"6F", x"6F", x"6E",
	x"6D", x"6D", x"6C", x"6C", x"6B", x"6C", x"6F", x"72", x"74", x"75", x"77", x"77",
	x"77", x"76", x"75", x"75", x"76", x"76", x"76", x"75", x"76", x"76", x"76", x"75",
	x"74", x"72", x"6E", x"6B", x"6A", x"6A", x"6A", x"6A", x"69", x"68", x"69", x"6B",
	x"6D", x"6F", x"6F", x"6E", x"6F", x"70", x"71", x"72", x"75", x"77", x"79", x"7A",
	x"7B", x"7B", x"7A", x"78", x"75", x"75", x"75", x"74", x"74", x"74", x"73", x"73",
	x"72", x"72", x"72", x"75", x"78", x"7A", x"7A", x"79", x"78", x"77", x"76", x"75",
	x"74", x"73", x"70", x"6E", x"6F", x"6E", x"6C", x"6B", x"6C", x"6C", x"6B", x"6A",
	x"68", x"66", x"64", x"61", x"60", x"5F", x"5E", x"5E", x"5F", x"61", x"64", x"68",
	x"6C", x"6F", x"71", x"72", x"72", x"72", x"73", x"72", x"70", x"6E", x"6D", x"6C",
	x"6A", x"67", x"65", x"64", x"65", x"67", x"69", x"69", x"68", x"65", x"61", x"5D",
	x"5A", x"59", x"57", x"56", x"55", x"54", x"50", x"4C", x"48", x"46", x"44", x"44",
	x"45", x"46", x"47", x"47", x"44", x"41", x"3F", x"3E", x"3D", x"3B", x"3A", x"38",
	x"37", x"38", x"38", x"38", x"39", x"38", x"36", x"35", x"34", x"35", x"37", x"3A",
	x"3C", x"3E", x"3E", x"3D", x"3A", x"36", x"31", x"2F", x"2E", x"2D", x"2C", x"2B",
	x"2A", x"29", x"26", x"23", x"21", x"1F", x"1D", x"1E", x"1F", x"1E", x"1C", x"19",
	x"18", x"19", x"1B", x"1B", x"1A", x"19", x"16", x"14", x"13", x"12", x"11", x"11",
	x"11", x"13", x"14", x"15", x"16", x"16", x"15", x"15", x"17", x"1A", x"1B", x"1B",
	x"1B", x"1B", x"1C", x"1C", x"1C", x"1D", x"1C", x"19", x"17", x"15", x"14", x"13",
	x"12", x"11", x"10", x"0F", x"10", x"12", x"12", x"10", x"0E", x"0B", x"09", x"07",
	x"05", x"03", x"03", x"04", x"03", x"00", x"FF", x"00", x"01", x"03", x"03", x"05",
	x"07", x"07", x"05", x"02", x"01", x"01", x"04", x"06", x"08", x"08", x"09", x"08",
	x"07", x"05", x"04", x"05", x"08", x"0A", x"0C", x"0D", x"0C", x"0C", x"0C", x"0B",
	x"0A", x"0B", x"09", x"07", x"04", x"02", x"01", x"02", x"03", x"06", x"09", x"0A",
	x"0B", x"0B", x"0B", x"0A", x"09", x"09", x"09", x"09", x"08", x"06", x"05", x"06",
	x"07", x"08", x"08", x"0A", x"0D", x"10", x"11", x"12", x"13", x"14", x"13", x"12",
	x"10", x"0F", x"0D", x"0D", x"0D", x"0C", x"0B", x"0B", x"0C", x"0C", x"0C", x"0D",
	x"0E", x"10", x"11", x"13", x"14", x"16", x"16", x"15", x"14", x"13", x"12", x"11",
	x"0F", x"0E", x"0E", x"0F", x"0E", x"0D", x"0B", x"09", x"08", x"07", x"05", x"04",
	x"04", x"05", x"08", x"08", x"07", x"07", x"07", x"07", x"08", x"08", x"06", x"04",
	x"02", x"00", x"FE", x"FD", x"FB", x"FB", x"FB", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FC", x"FD", x"FD", x"FC", x"FA", x"F9", x"F9", x"F8", x"F7", x"F6", x"F6", x"F6",
	x"F5", x"F5", x"F5", x"F8", x"F9", x"F9", x"FB", x"FC", x"FC", x"FC", x"FD", x"FD",
	x"FD", x"FE", x"00", x"00", x"00", x"FF", x"FC", x"F8", x"F5", x"F2", x"F0", x"ED",
	x"EC", x"EC", x"EC", x"EB", x"EC", x"ED", x"EE", x"EC", x"EA", x"E9", x"E7", x"E5",
	x"E4", x"E5", x"E5", x"E4", x"E4", x"E4", x"E3", x"E3", x"E2", x"E1", x"E1", x"E1",
	x"E1", x"E2", x"E1", x"E0", x"DF", x"DD", x"DB", x"D9", x"D8", x"D6", x"D6", x"D6",
	x"D6", x"D6", x"D5", x"D5", x"D4", x"D3", x"D2", x"D1", x"D1", x"D1", x"D2", x"D3",
	x"D4", x"D6", x"D8", x"DA", x"DA", x"DA", x"D9", x"D8", x"D6", x"D4", x"D0", x"CD",
	x"CB", x"CB", x"CC", x"CD", x"CD", x"CE", x"CF", x"D0", x"D1", x"D1", x"D1", x"D0",
	x"CF", x"CE", x"CD", x"CB", x"C9", x"C8", x"C9", x"C9", x"C8", x"C7", x"C7", x"C7",
	x"C8", x"C9", x"C9", x"C7", x"C5", x"C5", x"C5", x"C6", x"C6", x"C5", x"C3", x"C3",
	x"C3", x"C4", x"C5", x"C6", x"C7", x"C9", x"CB", x"CB", x"CA", x"C9", x"CA", x"C9",
	x"C8", x"C6", x"C3", x"C0", x"BD", x"BC", x"BD", x"C0", x"C2", x"C3", x"C4", x"C4",
	x"C3", x"C2", x"BF", x"BD", x"BB", x"B9", x"B7", x"B6", x"B7", x"B8", x"B8", x"B9",
	x"BB", x"BD", x"C1", x"C4", x"C5", x"C4", x"C5", x"C6", x"C5", x"C6", x"C7", x"C5",
	x"C3", x"C1", x"BF", x"BD", x"BA", x"B8", x"B7", x"B5", x"B3", x"B0", x"AD", x"AC",
	x"AB", x"AA", x"AC", x"AD", x"AE", x"B0", x"B1", x"B1", x"B2", x"B4", x"B6", x"B8",
	x"B9", x"B9", x"B9", x"B7", x"B7", x"B8", x"B9", x"BB", x"BB", x"BB", x"BB", x"BB",
	x"B9", x"B8", x"B7", x"B5", x"B3", x"B2", x"B1", x"B0", x"AF", x"AF", x"B0", x"B0",
	x"B1", x"B2", x"B3", x"B4", x"B5", x"B6", x"B6", x"B7", x"B8", x"B8", x"B8", x"BA",
	x"BC", x"BD", x"BE", x"BD", x"BC", x"BC", x"BE", x"BD", x"BA", x"B8", x"B7", x"B8",
	x"B8", x"B7", x"B6", x"B7", x"B8", x"B7", x"B7", x"B7", x"B9", x"BB", x"BC", x"BD",
	x"BE", x"BD", x"BE", x"BF", x"C0", x"C1", x"C2", x"C1", x"C0", x"C0", x"C1", x"C1",
	x"BF", x"BE", x"BE", x"BF", x"C1", x"C2", x"C3", x"C4", x"C6", x"C8", x"C8", x"C7",
	x"C6", x"C5", x"C6", x"C6", x"C7", x"C8", x"C9", x"CA", x"CA", x"CA", x"CC", x"CD",
	x"CD", x"CD", x"CE", x"D0", x"D2", x"D3", x"D4", x"D6", x"D6", x"D8", x"DB", x"DC",
	x"DB", x"DB", x"DA", x"DA", x"DB", x"DC", x"DB", x"D9", x"D8", x"D6", x"D5", x"D6",
	x"D6", x"D7", x"D9", x"DA", x"DB", x"DC", x"DE", x"DF", x"E0", x"DF", x"E1", x"E2",
	x"E3", x"E4", x"E4", x"E4", x"E4", x"E5", x"E5", x"E6", x"E7", x"EA", x"EC", x"ED",
	x"ED", x"EE", x"F0", x"F3", x"F6", x"F8", x"F9", x"F8", x"F8", x"F7", x"F5", x"F4",
	x"F2", x"F0", x"ED", x"EA", x"E8", x"E6", x"E5", x"E6", x"E7", x"E8", x"EA", x"ED",
	x"EF", x"F0", x"F2", x"F3", x"F3", x"F5", x"F6", x"F5", x"F4", x"F4", x"F5", x"F4",
	x"F3", x"F2", x"F3", x"F5", x"F6", x"F7", x"F8", x"F7", x"F6", x"F6", x"F7", x"F8",
	x"F7", x"F6", x"F5", x"F5", x"F4", x"F1", x"EE", x"ED", x"ED", x"EC", x"EB", x"EA",
	x"EB", x"EC", x"EC", x"EB", x"ED", x"EE", x"F1", x"F4", x"F6", x"F8", x"F9", x"F7",
	x"F6", x"F6", x"F5", x"F4", x"F3", x"F1", x"F0", x"EF", x"EE", x"EE", x"EE", x"EE",
	x"EE", x"EF", x"EF", x"F0", x"F2", x"F4", x"F5", x"F5", x"F4", x"F3", x"F2", x"F0",
	x"EF", x"ED", x"ED", x"EB", x"E8", x"E4", x"E1", x"E0", x"E0", x"E0", x"E1", x"E3",
	x"E4", x"E6", x"E7", x"E8", x"EA", x"EC", x"ED", x"EC", x"EC", x"ED", x"EF", x"F0",
	x"F1", x"F2", x"F3", x"F3", x"F2", x"F2", x"F1", x"F1", x"F2", x"F3", x"F3", x"F1",
	x"EE", x"EC", x"EC", x"EC", x"EA", x"E9", x"E9", x"E8", x"E6", x"E5", x"E3", x"E1",
	x"DE", x"DD", x"DE", x"DE", x"DE", x"E0", x"E2", x"E2", x"E5", x"E7", x"E9", x"EC",
	x"EE", x"F0", x"F1", x"F3", x"F4", x"F6", x"F9", x"FA", x"FA", x"F8", x"F6", x"F5",
	x"F5", x"F4", x"F2", x"F1", x"EF", x"EE", x"ED", x"ED", x"EC", x"ED", x"EF", x"F1",
	x"F2", x"F3", x"F4", x"F5", x"F6", x"F6", x"F7", x"F8", x"F8", x"F9", x"FA", x"F9",
	x"F8", x"F9", x"FA", x"FA", x"FB", x"FA", x"FA", x"FB", x"FB", x"FA", x"FA", x"FA",
	x"FC", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"FE", x"FD", x"FD", x"FE",
	x"00", x"02", x"02", x"03", x"04", x"07", x"0B", x"0D", x"0E", x"0D", x"0D", x"0D",
	x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0A", x"09", x"09", x"09", x"0A", x"0A",
	x"0A", x"0B", x"0B", x"0B", x"0C", x"0C", x"0D", x"0C", x"0C", x"0D", x"0E", x"10",
	x"12", x"15", x"17", x"18", x"1B", x"1E", x"1F", x"20", x"22", x"24", x"25", x"26",
	x"26", x"25", x"25", x"25", x"26", x"28", x"28", x"28", x"27", x"26", x"26", x"27",
	x"27", x"26", x"25", x"23", x"22", x"20", x"1E", x"1D", x"1E", x"1E", x"1E", x"1F",
	x"20", x"20", x"20", x"21", x"22", x"22", x"22", x"23", x"24", x"25", x"25", x"26",
	x"26", x"27", x"29", x"2A", x"2A", x"2A", x"29", x"28", x"27", x"28", x"29", x"29",
	x"29", x"2B", x"2C", x"2D", x"2D", x"2E", x"2F", x"2E", x"2C", x"2A", x"27", x"25",
	x"24", x"23", x"21", x"20", x"1F", x"1D", x"1D", x"1E", x"1E", x"20", x"22", x"22",
	x"23", x"25", x"25", x"25", x"23", x"22", x"22", x"22", x"22", x"22", x"23", x"24",
	x"25", x"25", x"26", x"26", x"27", x"26", x"25", x"23", x"20", x"1D", x"1C", x"1B",
	x"19", x"19", x"18", x"18", x"18", x"17", x"16", x"17", x"18", x"18", x"17", x"17",
	x"16", x"14", x"13", x"11", x"0F", x"0E", x"0D", x"0C", x"0B", x"09", x"08", x"06",
	x"04", x"03", x"02", x"00", x"FD", x"FC", x"FB", x"FA", x"F9", x"F9", x"FA", x"FB",
	x"FB", x"FC", x"FE", x"FF", x"FF", x"00", x"FF", x"FE", x"FC", x"FB", x"FA", x"F8",
	x"F7", x"F5", x"F3", x"F4", x"F5", x"F5", x"F5", x"F4", x"F5", x"F6", x"F7", x"F7",
	x"F7", x"F6", x"F5", x"F4", x"F4", x"F3", x"F1", x"EF", x"EE", x"ED", x"EB", x"E9",
	x"E9", x"E8", x"E8", x"E7", x"E7", x"E7", x"E7", x"E7", x"E7", x"E8", x"EA", x"EA",
	x"EB", x"EB", x"EB", x"EC", x"ED", x"ED", x"EE", x"EE", x"ED", x"EC", x"EB", x"EA",
	x"E9", x"E7", x"E6", x"E6", x"E6", x"E5", x"E5", x"E5", x"E4", x"E4", x"E6", x"E6",
	x"E6", x"E6", x"E7", x"E8", x"E9", x"E9", x"EA", x"EB", x"EC", x"ED", x"ED", x"EE",
	x"EE", x"EE", x"ED", x"EC", x"EC", x"EB", x"E9", x"E6", x"E5", x"E4", x"E4", x"E3",
	x"E1", x"E1", x"E2", x"E3", x"E5", x"E6", x"E6", x"E8", x"EB", x"EC", x"EC", x"ED",
	x"EE", x"EF", x"F0", x"EF", x"EF", x"EF", x"F0", x"F0", x"EF", x"ED", x"EC", x"EC",
	x"EC", x"EB", x"EC", x"ED", x"EE", x"F0", x"F1", x"F2", x"F4", x"F5", x"F5", x"F5",
	x"F4", x"F3", x"F3", x"F4", x"F4", x"F5", x"F5", x"F4", x"F4", x"F4", x"F5", x"F6",
	x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7",
	x"F8", x"F9", x"FA", x"FC", x"FD", x"FF", x"00", x"02", x"04", x"05", x"06", x"07",
	x"08", x"09", x"0B", x"0C", x"0E", x"0F", x"10", x"10", x"10", x"0F", x"0E", x"0D",
	x"0D", x"0C", x"0B", x"09", x"08", x"05", x"04", x"04", x"03", x"03", x"04", x"05",
	x"07", x"08", x"09", x"09", x"0A", x"0A", x"0B", x"0B", x"0B", x"0C", x"0C", x"0B",
	x"0B", x"0D", x"0F", x"10", x"10", x"0F", x"0F", x"0E", x"0E", x"10", x"11", x"10",
	x"0F", x"0E", x"0C", x"0A", x"09", x"09", x"0A", x"0A", x"0A", x"0B", x"0B", x"0B",
	x"0B", x"0C", x"0D", x"0E", x"0E", x"0F", x"10", x"11", x"13", x"14", x"15", x"17",
	x"19", x"19", x"18", x"16", x"15", x"15", x"14", x"13", x"12", x"11", x"0F", x"0F",
	x"0E", x"0F", x"10", x"11", x"11", x"10", x"11", x"12", x"12", x"13", x"13", x"14",
	x"15", x"15", x"15", x"15", x"16", x"16", x"16", x"16", x"18", x"1A", x"1A", x"1A",
	x"1A", x"1A", x"19", x"19", x"18", x"17", x"18", x"18", x"19", x"1A", x"1B", x"1A",
	x"1A", x"1B", x"1B", x"1B", x"1B", x"1B", x"1C", x"1B", x"1A", x"19", x"17", x"16",
	x"17", x"17", x"16", x"16", x"16", x"15", x"16", x"16", x"17", x"17", x"17", x"16",
	x"16", x"16", x"16", x"16", x"15", x"13", x"12", x"12", x"12", x"12", x"12", x"12",
	x"12", x"14", x"14", x"15", x"16", x"17", x"16", x"16", x"15", x"14", x"13", x"13",
	x"12", x"12", x"13", x"14", x"14", x"15", x"16", x"18", x"19", x"1A", x"1B", x"1C",
	x"1C", x"1D", x"1D", x"1C", x"1D", x"1C", x"1C", x"1C", x"1C", x"1B", x"1B", x"1C",
	x"1C", x"1B", x"19", x"19", x"19", x"1A", x"1A", x"1A", x"1A", x"1A", x"1A", x"1B",
	x"1B", x"1C", x"1D", x"1D", x"1C", x"1C", x"1B", x"1B", x"1B", x"1B", x"1C", x"1D",
	x"1E", x"1E", x"1E", x"1F", x"20", x"21", x"23", x"25", x"27", x"28", x"29", x"2B",
	x"2B", x"2B", x"2B", x"2C", x"2D", x"2C", x"2C", x"2B", x"2B", x"2A", x"29", x"29",
	x"29", x"28", x"27", x"27", x"26", x"25", x"24", x"23", x"22", x"23", x"23", x"22",
	x"22", x"21", x"21", x"21", x"21", x"22", x"23", x"24", x"24", x"24", x"25", x"25",
	x"25", x"25", x"25", x"25", x"25", x"24", x"24", x"24", x"24", x"24", x"24", x"23",
	x"23", x"23", x"24", x"23", x"23", x"22", x"23", x"23", x"22", x"21", x"21", x"20",
	x"1F", x"1F", x"1E", x"1E", x"20", x"20", x"20", x"1F", x"1E", x"1F", x"20", x"21",
	x"22", x"24", x"26", x"27", x"28", x"29", x"29", x"2A", x"29", x"29", x"2A", x"2C",
	x"2D", x"2E", x"2E", x"2F", x"31", x"32", x"32", x"31", x"31", x"32", x"32", x"32",
	x"32", x"32", x"33", x"33", x"33", x"34", x"33", x"33", x"32", x"31", x"31", x"31",
	x"31", x"30", x"2F", x"2F", x"2F", x"2F", x"2F", x"2F", x"2F", x"2F", x"2E", x"2F",
	x"30", x"31", x"32", x"32", x"31", x"30", x"31", x"31", x"31", x"32", x"32", x"33",
	x"34", x"34", x"35", x"35", x"35", x"35", x"37", x"38", x"39", x"39", x"3A", x"3B",
	x"3D", x"3D", x"3D", x"3D", x"3D", x"3D", x"3E", x"3E", x"3E", x"3E", x"3F", x"3F",
	x"3F", x"3F", x"3F", x"40", x"40", x"40", x"42", x"44", x"45", x"45", x"46", x"47",
	x"47", x"47", x"47", x"47", x"48", x"48", x"48", x"49", x"4A", x"4A", x"4A", x"4A",
	x"4B", x"4D", x"4D", x"4D", x"4E", x"4E", x"4D", x"4D", x"4D", x"4E", x"4F", x"4F",
	x"4E", x"4E", x"4D", x"4C", x"4D", x"4C", x"4C", x"4B", x"4A", x"49", x"49", x"49",
	x"48", x"47", x"47", x"48", x"48", x"4A", x"4B", x"4B", x"4B", x"4C", x"4D", x"4E",
	x"4F", x"50", x"51", x"51", x"51", x"52", x"52", x"51", x"51", x"50", x"4F", x"4F",
	x"4E", x"4D", x"4D", x"4C", x"4A", x"49", x"48", x"48", x"48", x"48", x"46", x"46",
	x"46", x"46", x"46", x"46", x"46", x"47", x"48", x"47", x"47", x"46", x"46", x"46",
	x"46", x"46", x"46", x"45", x"45", x"43", x"43", x"42", x"42", x"41", x"40", x"40",
	x"40", x"3F", x"3D", x"3B", x"3A", x"39", x"39", x"38", x"37", x"36", x"36", x"36",
	x"36", x"34", x"33", x"34", x"34", x"34", x"34", x"34", x"34", x"34", x"33", x"31",
	x"31", x"30", x"2F", x"2F", x"2F", x"2E", x"2E", x"2D", x"2C", x"2B", x"2B", x"2A",
	x"29", x"28", x"27", x"26", x"25", x"24", x"24", x"23", x"22", x"21", x"20", x"1F",
	x"1E", x"1E", x"1D", x"1C", x"1C", x"1C", x"1C", x"1C", x"1C", x"1B", x"1B", x"1A",
	x"1A", x"1A", x"1B", x"1B", x"1B", x"1A", x"18", x"16", x"15", x"14", x"13", x"11",
	x"0F", x"0E", x"0D", x"0C", x"0B", x"0A", x"09", x"09", x"09", x"08", x"07", x"07",
	x"06", x"06", x"06", x"05", x"04", x"04", x"02", x"01", x"FF", x"FE", x"FD", x"FC",
	x"FA", x"F9", x"F9", x"F9", x"F9", x"F8", x"F6", x"F4", x"F3", x"F3", x"F3", x"F3",
	x"F3", x"F3", x"F3", x"F3", x"F3", x"F4", x"F4", x"F4", x"F3", x"F2", x"F0", x"EF",
	x"EF", x"EE", x"ED", x"EC", x"EB", x"EB", x"EB", x"EA", x"EB", x"EB", x"EA", x"EA",
	x"E9", x"E9", x"E9", x"E8", x"E6", x"E4", x"E4", x"E4", x"E4", x"E4", x"E3", x"E3",
	x"E2", x"E1", x"E0", x"E0", x"E0", x"E0", x"E0", x"E0", x"DF", x"DE", x"DE", x"DF",
	x"DF", x"DE", x"DE", x"DE", x"DF", x"DE", x"DC", x"DB", x"D9", x"D8", x"D8", x"D8",
	x"D7", x"D7", x"D7", x"D6", x"D6", x"D5", x"D4", x"D5", x"D6", x"D6", x"D6", x"D6",
	x"D6", x"D7", x"D6", x"D5", x"D5", x"D4", x"D3", x"D2", x"D1", x"CE", x"CD", x"CC",
	x"CB", x"CB", x"CA", x"C9", x"C9", x"C8", x"C8", x"C9", x"CA", x"C9", x"C9", x"C9",
	x"C9", x"C8", x"C7", x"C7", x"C6", x"C6", x"C5", x"C4", x"C3", x"C2", x"C2", x"C1",
	x"C1", x"C0", x"C1", x"C1", x"C0", x"BF", x"BF", x"BF", x"BF", x"BF", x"BE", x"BE",
	x"BD", x"BD", x"BC", x"BB", x"BA", x"BA", x"B8", x"B8", x"B8", x"B8", x"B8", x"B9",
	x"B8", x"B8", x"B8", x"B7", x"B8", x"B8", x"B8", x"B8", x"B7", x"B8", x"B8", x"B7",
	x"B7", x"B6", x"B5", x"B4", x"B4", x"B4", x"B4", x"B3", x"B3", x"B3", x"B3", x"B3",
	x"B2", x"B2", x"B2", x"B2", x"B1", x"B0", x"B1", x"B1", x"B0", x"B0", x"B0", x"AF",
	x"AE", x"AE", x"AE", x"AE", x"AD", x"AC", x"AB", x"AA", x"AA", x"AB", x"AB", x"AA",
	x"AA", x"AA", x"AA", x"AA", x"AA", x"AA", x"A9", x"A9", x"A9", x"A9", x"AA", x"A9",
	x"A8", x"A7", x"A7", x"A6", x"A6", x"A5", x"A4", x"A4", x"A4", x"A4", x"A4", x"A3",
	x"A3", x"A3", x"A3", x"A3", x"A2", x"A2", x"A2", x"A3", x"A3", x"A3", x"A3", x"A3",
	x"A3", x"A2", x"A1", x"A1", x"A1", x"A0", x"A0", x"A0", x"A1", x"A0", x"9F", x"9F",
	x"9F", x"A0", x"A0", x"A0", x"A1", x"A3", x"A4", x"A4", x"A4", x"A4", x"A5", x"A6",
	x"A5", x"A4", x"A4", x"A5", x"A5", x"A5", x"A5", x"A4", x"A4", x"A5", x"A5", x"A6",
	x"A6", x"A6", x"A6", x"A8", x"A8", x"A9", x"A9", x"A9", x"A9", x"AA", x"A9", x"A8",
	x"A8", x"A8", x"A8", x"A7", x"A6", x"A6", x"A6", x"A7", x"A7", x"A7", x"A6", x"A6",
	x"A6", x"A6", x"A6", x"A7", x"A8", x"A9", x"AA", x"AB", x"AB", x"AB", x"AB", x"AB",
	x"AB", x"AB", x"AB", x"AB", x"AB", x"AB", x"AC", x"AC", x"AD", x"AD", x"AD", x"AD",
	x"AE", x"AE", x"AE", x"AE", x"AF", x"AF", x"AF", x"AF", x"B0", x"B1", x"B1", x"B2",
	x"B2", x"B2", x"B2", x"B3", x"B4", x"B3", x"B3", x"B2", x"B2", x"B2", x"B3", x"B3",
	x"B3", x"B4", x"B5", x"B6", x"B7", x"B8", x"B9", x"BA", x"BA", x"BA", x"BB", x"BB",
	x"BB", x"BC", x"BC", x"BC", x"BC", x"BC", x"BC", x"BD", x"BE", x"BF", x"C0", x"C1",
	x"C1", x"C2", x"C2", x"C2", x"C1", x"C1", x"C2", x"C2", x"C3", x"C3", x"C2", x"C2",
	x"C3", x"C3", x"C4", x"C5", x"C5", x"C5", x"C5", x"C5", x"C4", x"C3", x"C2", x"C2",
	x"C2", x"C2", x"C1", x"C1", x"C1", x"C1", x"C1", x"C1", x"C2", x"C3", x"C4", x"C3",
	x"C2", x"C1", x"C2", x"C4", x"C4", x"C5", x"C6", x"C6", x"C7", x"C7", x"C8", x"C9",
	x"CB", x"CC", x"CD", x"CE", x"CF", x"CF", x"D0", x"D0", x"D1", x"D1", x"D1", x"D2",
	x"D2", x"D1", x"D1", x"D2", x"D2", x"D3", x"D4", x"D5", x"D5", x"D4", x"D4", x"D3",
	x"D2", x"D2", x"D2", x"D2", x"D1", x"D1", x"D2", x"D1", x"D1", x"D1", x"D2", x"D2",
	x"D2", x"D2", x"D2", x"D3", x"D3", x"D3", x"D3", x"D3", x"D4", x"D5", x"D7", x"D7",
	x"D7", x"D8", x"DA", x"DA", x"DA", x"DA", x"DA", x"DB", x"DB", x"DB", x"DC", x"DC",
	x"DD", x"DD", x"DE", x"DF", x"E0", x"E0", x"E0", x"E1", x"E1", x"E1", x"E1", x"E1",
	x"E2", x"E2", x"E2", x"E2", x"E2", x"E2", x"E3", x"E3", x"E4", x"E4", x"E5", x"E5",
	x"E5", x"E5", x"E5", x"E4", x"E5", x"E7", x"E8", x"E8", x"E9", x"EA", x"EB", x"EB",
	x"EB", x"EA", x"EA", x"EA", x"EB", x"EB", x"EB", x"EB", x"EB", x"EB", x"EB", x"EB",
	x"EB", x"EB", x"EC", x"EB", x"EB", x"EB", x"EB", x"EC", x"EC", x"EC", x"EC", x"ED",
	x"ED", x"ED", x"EE", x"EF", x"F0", x"F1", x"F2", x"F2", x"F2", x"F2", x"F2", x"F3",
	x"F3", x"F2", x"F3", x"F4", x"F5", x"F5", x"F5", x"F5", x"F6", x"F7", x"F9", x"F9",
	x"FA", x"F9", x"F9", x"FA", x"FA", x"FA", x"FB", x"FC", x"FD", x"FD", x"FE", x"FE",
	x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"02", x"02", x"02", x"03", x"04",
	x"05", x"06", x"06", x"07", x"07", x"08", x"09", x"0A", x"09", x"09", x"0A", x"0B",
	x"0B", x"0C", x"0D", x"0D", x"0E", x"0F", x"0F", x"10", x"10", x"10", x"10", x"10",
	x"10", x"11", x"11", x"11", x"11", x"12", x"12", x"13", x"13", x"12", x"13", x"13",
	x"14", x"15", x"15", x"16", x"16", x"18", x"19", x"1A", x"1A", x"1B", x"1B", x"1D",
	x"1F", x"1F", x"20", x"20", x"20", x"21", x"21", x"21", x"21", x"21", x"21", x"21",
	x"21", x"22", x"23", x"23", x"24", x"24", x"24", x"24", x"24", x"25", x"24", x"24",
	x"25", x"25", x"26", x"27", x"26", x"27", x"27", x"27", x"28", x"28", x"28", x"28",
	x"29", x"29", x"29", x"29", x"28", x"28", x"29", x"29", x"28", x"28", x"27", x"27",
	x"27", x"27", x"27", x"27", x"27", x"27", x"27", x"27", x"27", x"27", x"27", x"27",
	x"27", x"27", x"28", x"29", x"29", x"29", x"29", x"28", x"28", x"28", x"28", x"28",
	x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"28", x"27", x"27", x"26", x"26",
	x"26", x"26", x"26", x"27", x"27", x"27", x"27", x"27", x"27", x"26", x"26", x"26",
	x"26", x"26", x"27", x"27", x"28", x"29", x"2A", x"2A", x"29", x"28", x"27", x"27",
	x"27", x"27", x"27", x"26", x"25", x"24", x"24", x"23", x"23", x"22", x"22", x"22",
	x"23", x"23", x"24", x"24", x"24", x"24", x"25", x"25", x"25", x"25", x"25", x"26",
	x"26", x"25", x"25", x"25", x"24", x"23", x"23", x"23", x"24", x"23", x"23", x"23",
	x"22", x"22", x"22", x"21", x"21", x"22", x"23", x"23", x"22", x"22", x"21", x"20",
	x"21", x"20", x"1F", x"1E", x"1D", x"1D", x"1D", x"1D", x"1D", x"1E", x"1E", x"1E",
	x"1F", x"1F", x"1F", x"20", x"1F", x"1F", x"1E", x"1E", x"1E", x"1E", x"1E", x"1E",
	x"1E", x"1E", x"1F", x"20", x"20", x"20", x"20", x"20", x"1F", x"20", x"21", x"21",
	x"22", x"22", x"23", x"23", x"23", x"22", x"22", x"22", x"21", x"20", x"20", x"1F",
	x"1F", x"1E", x"1D", x"1E", x"1E", x"1E", x"1E", x"1E", x"1D", x"1D", x"1E", x"1E",
	x"1F", x"1F", x"1F", x"1F", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"21",
	x"20", x"20", x"1F", x"1F", x"1E", x"1E", x"1D", x"1D", x"1D", x"1D", x"1D", x"1E",
	x"1E", x"1E", x"1E", x"1E", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F", x"1F",
	x"1E", x"1F", x"1F", x"1E", x"1E", x"1F", x"1F", x"1F", x"1E", x"1E", x"1E", x"1E",
	x"1F", x"1F", x"1F", x"1E", x"1E", x"1E", x"1E", x"1D", x"1D", x"1D", x"1D", x"1D",
	x"1E", x"1D", x"1D", x"1E", x"1E", x"1E", x"1E", x"1E", x"1F", x"1F", x"20", x"20",
	x"21", x"21", x"22", x"23", x"22", x"23", x"23", x"23", x"24", x"24", x"24", x"24",
	x"23", x"22", x"22", x"22", x"22", x"22", x"23", x"23", x"23", x"23", x"23", x"22",
	x"22", x"22", x"22", x"23", x"23", x"23", x"23", x"23", x"22", x"23", x"23", x"24",
	x"24", x"24", x"24", x"24", x"24", x"23", x"22", x"22", x"22", x"22", x"21", x"21",
	x"21", x"21", x"21", x"21", x"21", x"21", x"20", x"20", x"20", x"20", x"21", x"21",
	x"22", x"22", x"22", x"22", x"23", x"24", x"24", x"24", x"24", x"23", x"23", x"23",
	x"23", x"23", x"23", x"23", x"22", x"22", x"22", x"21", x"21", x"20", x"21", x"21",
	x"21", x"21", x"21", x"20", x"20", x"21", x"20", x"20", x"20", x"20", x"20", x"21",
	x"21", x"20", x"20", x"20", x"20", x"20", x"20", x"21", x"21", x"21", x"20", x"20",
	x"20", x"20", x"1F", x"1F", x"1F", x"1F", x"20", x"20", x"20", x"20", x"1F", x"20",
	x"20", x"1F", x"1F", x"1F", x"1F", x"20", x"20", x"20", x"20", x"20", x"1F", x"20",
	x"20", x"20", x"20", x"20", x"1F", x"1F", x"20", x"1F", x"1F", x"1F", x"1E", x"1E",
	x"1F", x"1F", x"1E", x"1E", x"1E", x"1E", x"1F", x"1F", x"1F", x"1F", x"1E", x"1D",
	x"1C", x"1C", x"1B", x"1B", x"1A", x"1A", x"1A", x"1A", x"19", x"19", x"19", x"19",
	x"19", x"19", x"18", x"18", x"18", x"18", x"19", x"19", x"19", x"1A", x"1B", x"1B",
	x"1B", x"1B", x"1A", x"1B", x"1C", x"1B", x"1B", x"1C", x"1B", x"1B", x"1B", x"1B",
	x"1A", x"1B", x"1B", x"1A", x"1A", x"1A", x"1A", x"1A", x"1A", x"1A", x"1A", x"1A",
	x"1A", x"1A", x"1A", x"19", x"19", x"1A", x"19", x"19", x"19", x"19", x"19", x"19",
	x"19", x"19", x"19", x"19", x"19", x"19", x"19", x"19", x"18", x"18", x"18", x"18",
	x"18", x"17", x"17", x"16", x"16", x"16", x"16", x"15", x"15", x"14", x"14", x"14",
	x"14", x"13", x"13", x"13", x"12", x"12", x"12", x"12", x"13", x"13", x"13", x"13",
	x"13", x"12", x"12", x"11", x"11", x"11", x"11", x"10", x"10", x"10", x"10", x"0F",
	x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"10", x"0F", x"0F",
	x"0F", x"0E", x"0E", x"0F", x"0E", x"0D", x"0D", x"0C", x"0C", x"0B", x"0A", x"09",
	x"09", x"09", x"09", x"08", x"07", x"06", x"05", x"05", x"05", x"05", x"05", x"04",
	x"04", x"04", x"03", x"03", x"03", x"03", x"03", x"03", x"04", x"04", x"04", x"04",
	x"03", x"04", x"03", x"03", x"03", x"03", x"02", x"02", x"02", x"01", x"00", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE",
	x"FD", x"FD", x"FD", x"FC", x"FC", x"FC", x"FB", x"FB", x"FB", x"FA", x"FA", x"F9",
	x"F8", x"F8", x"F7", x"F6", x"F6", x"F7", x"F6", x"F6", x"F6", x"F5", x"F5", x"F6",
	x"F6", x"F6", x"F6", x"F6", x"F5", x"F6", x"F5", x"F5", x"F5", x"F4", x"F2", x"F2",
	x"F2", x"F2", x"F2", x"F1", x"F1", x"F1", x"F1", x"F1", x"F0", x"F0", x"F0", x"F0",
	x"F1", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"EF", x"EF", x"EF", x"EF", x"EF",
	x"EF", x"EF", x"EF", x"EF", x"EE", x"EE", x"EF", x"EE", x"EE", x"EE", x"EE", x"EE",
	x"EE", x"EE", x"EE", x"EE", x"EF", x"EF", x"EF", x"EE", x"ED", x"ED", x"ED", x"EE",
	x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"ED", x"ED", x"ED", x"ED",
	x"ED", x"EE", x"EE", x"ED", x"ED", x"ED", x"ED", x"ED", x"EC", x"EC", x"EC", x"EC",
	x"EC", x"EC", x"EC", x"EB", x"EB", x"EB", x"EB", x"EC", x"EC", x"EC", x"EC", x"EC",
	x"EC", x"EB", x"EB", x"EB", x"EB", x"EB", x"EB", x"EC", x"EC", x"EC", x"EC", x"EC",
	x"EC", x"ED", x"ED", x"EC", x"EC", x"EC", x"EC", x"EC", x"ED", x"ED", x"ED", x"ED",
	x"ED", x"EE", x"EE", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"F0",
	x"F0", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F2", x"F2", x"F1", x"F0", x"F0",
	x"F1", x"F1", x"F1", x"F0", x"F0", x"F0", x"F1", x"F1", x"F1", x"F1", x"F0", x"F0",
	x"F1", x"F0", x"F0", x"F0", x"F0", x"F0", x"F1", x"F0", x"F0", x"F0", x"F0", x"F0",
	x"F1", x"F1", x"F0", x"F1", x"F1", x"F2", x"F2", x"F2", x"F2", x"F3", x"F3", x"F3",
	x"F3", x"F3", x"F3", x"F3", x"F4", x"F4", x"F4", x"F4", x"F4", x"F4", x"F4", x"F3",
	x"F4", x"F4", x"F4", x"F4", x"F4", x"F4", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3",
	x"F3", x"F3", x"F2", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F4", x"F4",
	x"F4", x"F4", x"F3", x"F3", x"F4", x"F3", x"F3", x"F3", x"F3", x"F3", x"F2", x"F2",
	x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F2", x"F3",
	x"F3", x"F4", x"F4", x"F4", x"F5", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6",
	x"F6", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F4", x"F4", x"F3", x"F3",
	x"F3", x"F3", x"F3", x"F2", x"F2", x"F2", x"F3", x"F2", x"F2", x"F2", x"F2", x"F2",
	x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F2", x"F2", x"F2", x"F2", x"F2",
	x"F2", x"F2", x"F2", x"F2", x"F1", x"F1", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2",
	x"F2", x"F2", x"F2", x"F2", x"F2", x"F3", x"F3", x"F3", x"F2", x"F2", x"F2", x"F2",
	x"F2", x"F2", x"F2", x"F3", x"F3", x"F3", x"F2", x"F2", x"F2", x"F2", x"F3", x"F2",
	x"F2", x"F2", x"F2", x"F1", x"F1", x"F1", x"F1", x"F2", x"F1", x"F1", x"F1", x"F1",
	x"F1", x"F1", x"F1", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0",
	x"F0", x"F0", x"F0", x"F0", x"F0", x"F1", x"F1", x"F1", x"F2", x"F2", x"F2", x"F2",
	x"F2", x"F2", x"F2", x"F2", x"F2", x"F3", x"F3", x"F3", x"F3", x"F2", x"F2", x"F3",
	x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F2", x"F2", x"F1", x"F2",
	x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F1", x"F1", x"F1", x"F1", x"F2",
	x"F2", x"F3", x"F3", x"F3", x"F2", x"F2", x"F2", x"F2", x"F2", x"F1", x"F1", x"F1",
	x"F2", x"F2", x"F2", x"F2", x"F2", x"F3", x"F3", x"F3", x"F3", x"F4", x"F4", x"F4",
	x"F3", x"F4", x"F4", x"F4", x"F4", x"F4", x"F4", x"F4", x"F4", x"F4", x"F3", x"F3",
	x"F3", x"F3", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2",
	x"F2", x"F3", x"F2", x"F2", x"F2", x"F2", x"F3", x"F3", x"F2", x"F2", x"F2", x"F2",
	x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F3", x"F3", x"F3", x"F3",
	x"F2", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F2", x"F2", x"F2", x"F2",
	x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F1", x"F2", x"F2", x"F1", x"F1", x"F1",
	x"F1", x"F1", x"F2", x"F2", x"F2", x"F2", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1",
	x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0",
	x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"EF", x"F0", x"EF", x"EF", x"EF",
	x"F0", x"EF", x"F0", x"F0", x"EF", x"EF", x"EF", x"EE", x"EF", x"EF", x"EE", x"EE",
	x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EF", x"EE", x"EE",
	x"EE", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"F0", x"F0", x"EF",
	x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"EF", x"F0", x"F0", x"F0",
	x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F1", x"F1", x"F0",
	x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F0", x"F1", x"F1", x"F1", x"F2", x"F2",
	x"F2", x"F2", x"F2", x"F2", x"F2", x"F3", x"F3", x"F4", x"F4", x"F4", x"F4", x"F4",
	x"F4", x"F5", x"F5", x"F5", x"F5", x"F5", x"F4", x"F4", x"F4", x"F4", x"F3", x"F3",
	x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F3", x"F4", x"F4",
	x"F4", x"F5", x"F5", x"F4", x"F4", x"F5", x"F5", x"F5", x"F6", x"F6", x"F6", x"F7",
	x"F7", x"F7", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F9", x"F9",
	x"FA", x"F9", x"FA", x"FA", x"F9", x"F9", x"FA", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FB", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FD", x"FD", x"FC", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"01", x"01", x"01", x"02", x"02", x"02", x"03", x"02", x"02", x"03",
	x"03", x"03", x"03", x"03", x"04", x"04", x"04", x"04", x"05", x"05", x"05", x"05",
	x"04", x"04", x"04", x"04", x"04", x"05", x"05", x"04", x"05", x"04", x"04", x"05",
	x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05",
	x"05", x"05", x"05", x"06", x"06", x"06", x"06", x"06", x"06", x"07", x"06", x"06",
	x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"05",
	x"05", x"05", x"05", x"05", x"05", x"05", x"06", x"06", x"06", x"06", x"06", x"06",
	x"07", x"07", x"07", x"08", x"08", x"08", x"08", x"08", x"09", x"09", x"0A", x"0A",
	x"0A", x"0A", x"0A", x"0B", x"0B", x"0B", x"0A", x"0B", x"0B", x"0B", x"0B", x"0B",
	x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0B", x"0A", x"0A", x"0A", x"0B",
	x"0B", x"0B", x"0B", x"0B", x"0B", x"0A", x"0A", x"0A", x"0A", x"0B", x"0B", x"0B",
	x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0A", x"0B", x"0B", x"0B", x"0B", x"0C",
	x"0B", x"0C", x"0C", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0C", x"0C", x"0C",
	x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0D", x"0D", x"0D", x"0D", x"0D",
	x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0C",
	x"0C", x"0C", x"0C", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D",
	x"0D", x"0D", x"0D", x"0E", x"0E", x"0E", x"0E", x"0E", x"0E", x"0E", x"0E", x"0F",
	x"0F", x"0E", x"0E", x"0F", x"0F", x"0F", x"0F", x"0E", x"0E", x"0E", x"0E", x"0E",
	x"0E", x"0E", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0D", x"0C", x"0C", x"0C",
	x"0C", x"0C", x"0B", x"0C", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B", x"0B",
	x"0A", x"0A", x"0B", x"0B", x"0B", x"0B", x"0A", x"0B", x"0A", x"0A", x"0A", x"0A",
	x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A",
	x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", x"09", x"09", x"09", x"0A", x"0A", x"0A",
	x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09",
	x"09", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08",
	x"08", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07",
	x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07",
	x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"06", x"06", x"06", x"06", x"06",
	x"06", x"06", x"06", x"07", x"07", x"06", x"07", x"06", x"06", x"06", x"06", x"06",
	x"06", x"06", x"06", x"06", x"06", x"05", x"05", x"05", x"05", x"05", x"05", x"05",
	x"06", x"06", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"06",
	x"06", x"07", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06",
	x"06", x"06", x"06", x"05", x"06", x"06", x"05", x"05", x"05", x"04", x"04", x"04",
	x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"03", x"04", x"03",
	x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"02", x"03", x"02", x"02", x"02",
	x"02", x"02", x"02", x"02", x"02", x"03", x"02", x"02", x"02", x"02", x"02", x"02",
	x"03", x"03", x"03", x"02", x"02", x"02", x"02", x"01", x"01", x"02", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FD", x"FC", x"FC", x"FC", x"FC", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"FA", x"FA", x"FA", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"F9", x"F8", x"F8", x"F8", x"F9", x"F9", x"F9", x"F8",
	x"F8", x"F8", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"F6", x"F5", x"F5", x"F6",
	x"F5", x"F6", x"F6", x"F6", x"F6", x"F6", x"F5", x"F5", x"F6", x"F5", x"F6", x"F6",
	x"F6", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F6", x"F6", x"F6", x"F6",
	x"F5", x"F5", x"F6", x"F6", x"F5", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6",
	x"F6", x"F6", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5",
	x"F5", x"F5", x"F6", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5",
	x"F6", x"F6", x"F6", x"F6", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7",
	x"F8", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F8", x"F8", x"F8",
	x"F8", x"F8", x"F8", x"F8", x"F9", x"F8", x"F8", x"F8", x"F8", x"F8", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"F9", x"F8", x"F8", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"F9", x"F9", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FB",
	x"FB", x"FA", x"FA", x"FA", x"FA", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FA", x"FA", x"FA", x"FA", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02",
	x"02", x"02", x"02", x"02", x"02", x"02", x"01", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD",
	x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FC", x"FC", x"FC", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"01", x"01", x"01", x"00", x"01", x"01", x"01", x"01", x"01", x"00",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"02", x"01", x"01",
	x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"03", x"03", x"03",
	x"03", x"03", x"03", x"03", x"03", x"04", x"03", x"04", x"04", x"04", x"05", x"05",
	x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"06", x"06",
	x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"07", x"07",
	x"06", x"06", x"06", x"06", x"06", x"07", x"07", x"07", x"07", x"07", x"07", x"07",
	x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07",
	x"07", x"07", x"07", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06",
	x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"05", x"05", x"05", x"05", x"05",
	x"06", x"05", x"05", x"05", x"05", x"05", x"06", x"05", x"05", x"06", x"05", x"05",
	x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"06", x"05",
	x"05", x"05", x"05", x"06", x"06", x"05", x"05", x"05", x"05", x"05", x"06", x"05",
	x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"04", x"04", x"04", x"04",
	x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"03", x"03", x"03", x"03",
	x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"02", x"02",
	x"02", x"01", x"02", x"02", x"02", x"02", x"02", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FC", x"FD", x"FD", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F8",
	x"F8", x"F8", x"F8", x"F8", x"F8", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7",
	x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7",
	x"F7", x"F7", x"F7", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6",
	x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6",
	x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F7",
	x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F8", x"F7", x"F7", x"F7",
	x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F8",
	x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8",
	x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"FA", x"FA", x"FA", x"FA", x"FA", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"01", x"01", x"01", x"01", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02",
	x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02",
	x"02", x"02", x"03", x"02", x"02", x"03", x"03", x"03", x"03", x"03", x"03", x"04",
	x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"05", x"05", x"05", x"05",
	x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"06", x"06", x"06", x"06",
	x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06",
	x"06", x"06", x"06", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05",
	x"05", x"05", x"04", x"05", x"05", x"05", x"05", x"05", x"04", x"04", x"04", x"05",
	x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05",
	x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05",
	x"05", x"05", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"03", x"04", x"04",
	x"04", x"04", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03",
	x"03", x"03", x"03", x"03", x"03", x"03", x"02", x"02", x"03", x"02", x"02", x"02",
	x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02",
	x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"01", x"01", x"02",
	x"02", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"01", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD",
	x"FE", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FC", x"FD", x"FC", x"FC", x"FD", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FB", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FA", x"FB",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"F9", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"F9", x"F9", x"FA", x"FA", x"FA", x"FA", x"FA", x"F9", x"FA", x"FA", x"F9",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"F9", x"F9", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"FA", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"FA", x"FA", x"F9", x"F9", x"F9", x"FA", x"FA", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"FA", x"FA", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"02", x"02", x"02",
	x"02", x"02", x"02", x"02", x"02", x"02", x"03", x"03", x"03", x"03", x"03", x"03",
	x"03", x"03", x"03", x"03", x"04", x"03", x"04", x"04", x"04", x"04", x"04", x"04",
	x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"05",
	x"05", x"05", x"04", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05",
	x"05", x"05", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"05", x"06", x"06",
	x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"06",
	x"06", x"06", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07",
	x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07",
	x"08", x"07", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"09", x"09", x"09",
	x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09",
	x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09",
	x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09", x"09",
	x"09", x"09", x"09", x"09", x"09", x"08", x"08", x"08", x"08", x"08", x"08", x"08",
	x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"07", x"08", x"08",
	x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08",
	x"07", x"08", x"08", x"07", x"07", x"07", x"07", x"08", x"08", x"08", x"08", x"08",
	x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08",
	x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"07", x"07",
	x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07",
	x"07", x"07", x"07", x"07", x"06", x"06", x"07", x"06", x"06", x"06", x"06", x"06",
	x"06", x"06", x"06", x"06", x"06", x"06", x"06", x"05", x"05", x"05", x"05", x"05",
	x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05", x"05",
	x"05", x"05", x"05", x"05", x"05", x"04", x"04", x"04", x"04", x"04", x"04", x"04",
	x"04", x"04", x"04", x"04", x"04", x"04", x"03", x"04", x"03", x"03", x"03", x"03",
	x"03", x"03", x"03", x"02", x"03", x"03", x"02", x"03", x"02", x"02", x"02", x"02",
	x"02", x"02", x"02", x"02", x"02", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FA", x"FB", x"FB", x"FB", x"FB", x"FB", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"F9", x"F9", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"F9", x"FA", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F9",
	x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8",
	x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8",
	x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8",
	x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FB", x"FB", x"FB", x"FB", x"FB", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FB", x"FA", x"FA", x"FB",
	x"FA", x"FA", x"FB", x"FA", x"FA", x"FB", x"FA", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FA", x"FB", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"F9", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FB", x"FB", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FA", x"FA", x"FB", x"FA", x"FA", x"FB", x"FA", x"FA", x"FA", x"FA", x"FA", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FC", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FC", x"FB", x"FC", x"FB", x"FB", x"FB", x"FB", x"FB", x"FC", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FE",
	x"FE", x"FE", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"02", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"02", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"02", x"02", x"01", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02",
	x"02", x"01", x"02", x"01", x"01", x"02", x"02", x"02", x"02", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"01",
	x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"01", x"00",
	x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00",
	x"01", x"01", x"00", x"00", x"01", x"00", x"00", x"01", x"00", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"02",
	x"01", x"01", x"02", x"01", x"01", x"02", x"02", x"01", x"02", x"01", x"01", x"02",
	x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02",
	x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"03", x"02", x"02",
	x"03", x"03", x"02", x"02", x"02", x"02", x"03", x"03", x"03", x"03", x"03", x"02",
	x"03", x"02", x"02", x"03", x"03", x"02", x"03", x"03", x"02", x"03", x"03", x"03",
	x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"02", x"03", x"03", x"03",
	x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03",
	x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03",
	x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03",
	x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03",
	x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03",
	x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"02", x"03", x"03", x"02", x"03",
	x"03", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02",
	x"02", x"02", x"01", x"01", x"01", x"02", x"02", x"01", x"01", x"02", x"02", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FD", x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FB", x"FB", x"FC", x"FB", x"FB",
	x"FC", x"FC", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FC",
	x"FC", x"FB", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"01", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"01", x"01", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"01", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"01", x"01",
	x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"02", x"01", x"02", x"02", x"02", x"02",
	x"02", x"02", x"01", x"02", x"02", x"01", x"02", x"02", x"02", x"02", x"02", x"02",
	x"02", x"02", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00"	
);

signal cnt_out: integer := 0;	
signal play_sound: std_logic := '0';
constant cnt_max: integer := 9557;
--signal out_signal: signed(7 downto 0) := x"00";

begin

process (CLK)
begin
    if rising_edge(CLK) then
        if RST = '1' then
            play_sound <= '0';
        elsif PLAY = '1' then
            play_sound <= '1';
        elsif PLAY = '0' and cnt_out = cnt_max then
            play_sound <= '0';
        end if;
    end if;
end process;

	
-- 12bit counter
process (CLK)
begin     
    if rising_edge(CLK) then
        if RST = '1' then
            cnt_out <= 0;
        elsif CE = '1' and play_sound = '1' then
            cnt_out <= cnt_out + 1;       
        end if;
        if cnt_out = cnt_max then
            cnt_out <= 0;            
        end if;        
    end if;
end process;

--SAMPLE_OUT <= kick_sound(conv_integer(cnt_out));
process (CLK) 
begin
    if rising_edge(CLK) then
        if RST = '1' then
            KICK_SAMP_O <= x"00";
        elsif CE = '1' then
            KICK_SAMP_O <= kick_sound(cnt_out);
        end if;
    end if;    
end process;

end Behavioral;
