----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 25.12.2018 17:39:59
-- Design Name: 
-- Module Name: Tom1 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Tom1 is
    Port ( CLK : in STD_LOGIC;
           CE : in STD_LOGIC;
           RST : in STD_LOGIC;
           PLAY : in STD_LOGIC;
           SAMPLE_OUT : out signed(7 downto 0)
           );
end Tom1;

architecture Behavioral of Tom1 is

type memory is array (0 to 8959) of signed(7 downto 0);
constant tom1_sound: memory := (
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"01", x"00", x"01", x"00",
	x"01", x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"01", x"00", x"01",
	x"00", x"01", x"00", x"01", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FC", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD", x"FC", x"FC", x"FC", x"FB", x"FC",
	x"FB", x"FC", x"FB", x"FB", x"FC", x"FA", x"FC", x"FB", x"FA", x"FB", x"FA", x"FB",
	x"FB", x"FB", x"FA", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FC", x"FB", x"FB",
	x"FC", x"FC", x"FB", x"FD", x"FB", x"FD", x"FB", x"FD", x"FB", x"FE", x"FC", x"FE",
	x"FC", x"FF", x"FC", x"FF", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"00", x"FB",
	x"03", x"EC", x"BC", x"AB", x"A5", x"9B", x"AB", x"98", x"C2", x"9B", x"BB", x"FE",
	x"E5", x"FD", x"EE", x"40", x"55", x"45", x"50", x"45", x"3F", x"3D", x"3D", x"0D",
	x"27", x"23", x"1B", x"0A", x"02", x"2D", x"E4", x"39", x"28", x"DF", x"10", x"03",
	x"20", x"2E", x"24", x"20", x"17", x"10", x"19", x"00", x"F3", x"14", x"00", x"FF",
	x"03", x"D6", x"CF", x"C7", x"BD", x"BE", x"BF", x"B4", x"C2", x"BB", x"BB", x"BD",
	x"B1", x"B6", x"BF", x"BA", x"BE", x"CA", x"C9", x"E4", x"EE", x"08", x"00", x"18",
	x"36", x"4D", x"5E", x"5F", x"66", x"43", x"62", x"52", x"39", x"42", x"30", x"29",
	x"1F", x"38", x"23", x"12", x"0A", x"0E", x"FA", x"EC", x"DE", x"C5", x"E1", x"D5",
	x"E6", x"D2", x"C7", x"CE", x"D2", x"E3", x"DB", x"E1", x"EE", x"02", x"F7", x"EE",
	x"F8", x"07", x"FE", x"DC", x"DE", x"E9", x"EE", x"E6", x"DA", x"DB", x"E7", x"E0",
	x"D5", x"EE", x"F3", x"FD", x"FB", x"00", x"16", x"29", x"37", x"2C", x"40", x"44",
	x"3A", x"3B", x"41", x"51", x"47", x"4D", x"46", x"41", x"39", x"2F", x"27", x"06",
	x"13", x"E7", x"D3", x"C4", x"B0", x"B9", x"AD", x"B8", x"AB", x"B7", x"C4", x"BE",
	x"B9", x"B3", x"C0", x"C4", x"C2", x"D2", x"D7", x"FF", x"1C", x"22", x"2D", x"2C",
	x"3A", x"33", x"40", x"45", x"41", x"37", x"37", x"29", x"23", x"2B", x"1C", x"14",
	x"10", x"0C", x"01", x"FA", x"F4", x"FF", x"0D", x"08", x"FE", x"09", x"0D", x"10",
	x"0B", x"0D", x"FE", x"09", x"0E", x"FB", x"0A", x"05", x"EF", x"E0", x"DD", x"DA",
	x"D7", x"CE", x"CC", x"C3", x"C5", x"BF", x"BD", x"BE", x"BD", x"C5", x"CE", x"DB",
	x"D4", x"E1", x"E9", x"F1", x"07", x"1D", x"33", x"35", x"4A", x"4D", x"4E", x"58",
	x"50", x"45", x"3B", x"43", x"3E", x"35", x"33", x"22", x"23", x"13", x"02", x"ED",
	x"DB", x"D7", x"CC", x"CA", x"C6", x"C7", x"CD", x"D3", x"CE", x"C9", x"CE", x"C8",
	x"DA", x"E9", x"DE", x"E8", x"EC", x"F3", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE",
	x"F9", x"ED", x"EE", x"F5", x"02", x"07", x"0A", x"08", x"08", x"09", x"10", x"15",
	x"1C", x"26", x"27", x"30", x"2F", x"35", x"31", x"35", x"37", x"30", x"31", x"1F",
	x"13", x"1F", x"1B", x"1A", x"0A", x"FA", x"F2", x"E2", x"DC", x"CB", x"C7", x"CA",
	x"CE", x"CE", x"CE", x"CD", x"C7", x"C9", x"D0", x"D7", x"CB", x"CB", x"D2", x"DE",
	x"ED", x"F2", x"FC", x"0B", x"19", x"1E", x"1D", x"13", x"21", x"2C", x"2E", x"32",
	x"31", x"2F", x"2C", x"30", x"2C", x"2E", x"2A", x"2A", x"29", x"20", x"14", x"0A",
	x"04", x"03", x"05", x"03", x"07", x"06", x"00", x"F8", x"EC", x"E6", x"E0", x"D8",
	x"D1", x"D3", x"DB", x"D7", x"DB", x"CE", x"D0", x"D5", x"D9", x"D4", x"CA", x"CE",
	x"D4", x"E2", x"E5", x"EB", x"EF", x"FD", x"0B", x"0A", x"11", x"1C", x"27", x"2F",
	x"2A", x"22", x"26", x"27", x"30", x"33", x"33", x"2D", x"29", x"26", x"1B", x"10",
	x"15", x"16", x"21", x"1F", x"19", x"16", x"0D", x"04", x"FC", x"F7", x"EB", x"E3",
	x"D7", x"D3", x"D2", x"D3", x"D2", x"CB", x"CD", x"C7", x"C8", x"C0", x"C2", x"C6",
	x"CC", x"DA", x"E0", x"EB", x"EB", x"F1", x"FB", x"04", x"0A", x"10", x"1B", x"25",
	x"2A", x"29", x"30", x"33", x"2F", x"2B", x"24", x"20", x"25", x"2B", x"34", x"35",
	x"33", x"2C", x"21", x"1D", x"12", x"09", x"FB", x"F5", x"F3", x"F2", x"EA", x"E4",
	x"F0", x"EC", x"F3", x"E9", x"EE", x"E5", x"E1", x"E2", x"D8", x"D7", x"D1", x"D0",
	x"D1", x"D0", x"D1", x"D1", x"D2", x"DB", x"DB", x"E0", x"E5", x"EB", x"FA", x"FB",
	x"03", x"09", x"1B", x"22", x"2E", x"2F", x"2E", x"2C", x"2B", x"2C", x"2E", x"32",
	x"2E", x"35", x"32", x"36", x"36", x"30", x"27", x"18", x"0D", x"04", x"FC", x"F5",
	x"F7", x"ED", x"E0", x"DE", x"DF", x"D0", x"CC", x"CF", x"CE", x"CF", x"D0", x"CF",
	x"D5", x"E3", x"E5", x"E6", x"E2", x"E2", x"E6", x"EA", x"EF", x"F6", x"F7", x"F3",
	x"FB", x"FC", x"FE", x"FE", x"06", x"08", x"0D", x"10", x"1C", x"28", x"2B", x"2A",
	x"2E", x"30", x"2C", x"28", x"2A", x"32", x"32", x"33", x"28", x"20", x"18", x"11",
	x"13", x"09", x"02", x"FC", x"F9", x"F2", x"E6", x"DE", x"DD", x"D6", x"D1", x"D0",
	x"D0", x"CA", x"CC", x"CB", x"CD", x"CD", x"D2", x"DB", x"E2", x"E6", x"E5", x"EB",
	x"EB", x"F3", x"F2", x"FC", x"02", x"0B", x"12", x"16", x"1F", x"21", x"28", x"2A",
	x"33", x"31", x"30", x"28", x"23", x"26", x"20", x"17", x"12", x"11", x"0E", x"13",
	x"1A", x"15", x"1C", x"15", x"0E", x"05", x"FE", x"FD", x"F5", x"F4", x"F1", x"EB",
	x"E8", x"E5", x"DE", x"D7", x"D1", x"C9", x"C6", x"C6", x"C2", x"C6", x"C9", x"D0",
	x"D9", x"DE", x"E6", x"EA", x"F6", x"FB", x"FF", x"07", x"0B", x"13", x"1B", x"1B",
	x"22", x"25", x"2C", x"35", x"33", x"32", x"30", x"2E", x"2A", x"27", x"22", x"20",
	x"1B", x"1B", x"15", x"0B", x"08", x"FF", x"FC", x"FA", x"F5", x"FD", x"FA", x"F1",
	x"F0", x"EB", x"E2", x"DF", x"DE", x"E1", x"E3", x"E4", x"E5", x"E4", x"E3", x"E1",
	x"DE", x"DF", x"DA", x"E0", x"E2", x"E1", x"E3", x"E3", x"EF", x"EF", x"F1", x"F8",
	x"FD", x"FF", x"06", x"0D", x"15", x"1F", x"27", x"2E", x"34", x"39", x"3C", x"3B",
	x"38", x"33", x"30", x"2F", x"31", x"27", x"1A", x"17", x"0D", x"01", x"FB", x"F2",
	x"EE", x"E7", x"E0", x"DD", x"DA", x"DA", x"D9", x"D9", x"DC", x"DC", x"DD", x"DD",
	x"DD", x"E1", x"E3", x"E2", x"E2", x"E4", x"EA", x"E6", x"E9", x"F0", x"F6", x"FE",
	x"FC", x"00", x"01", x"05", x"09", x"0E", x"0E", x"15", x"16", x"1C", x"1C", x"18",
	x"1B", x"19", x"1F", x"20", x"1F", x"1F", x"1D", x"22", x"20", x"1D", x"21", x"1D",
	x"1F", x"18", x"18", x"11", x"09", x"01", x"FB", x"F0", x"E4", x"E0", x"D7", x"D6",
	x"D0", x"D2", x"CE", x"D1", x"D3", x"D0", x"D4", x"D6", x"D9", x"DD", x"E4", x"EA",
	x"EC", x"F3", x"F6", x"F9", x"FF", x"02", x"05", x"0B", x"11", x"12", x"17", x"19",
	x"18", x"1E", x"1F", x"20", x"23", x"28", x"25", x"25", x"24", x"24", x"20", x"1C",
	x"16", x"13", x"0E", x"0E", x"0A", x"03", x"00", x"01", x"FB", x"FA", x"FA", x"F2",
	x"ED", x"EE", x"E5", x"E3", x"E2", x"E6", x"E4", x"DF", x"DB", x"DD", x"DD", x"D7",
	x"D7", x"D7", x"D8", x"DF", x"E2", x"E6", x"E9", x"F0", x"F9", x"FA", x"04", x"09",
	x"0D", x"12", x"18", x"1B", x"1D", x"22", x"27", x"25", x"26", x"27", x"28", x"2C",
	x"2A", x"25", x"1E", x"18", x"11", x"10", x"0E", x"0B", x"06", x"04", x"00", x"FF",
	x"FB", x"F4", x"F4", x"F1", x"F1", x"EF", x"EE", x"ED", x"E7", x"E2", x"DC", x"D8",
	x"DA", x"D8", x"DB", x"D9", x"DA", x"DD", x"DE", x"E3", x"EB", x"EC", x"EF", x"F5",
	x"F7", x"FE", x"FF", x"04", x"0E", x"0E", x"11", x"1B", x"1F", x"1F", x"24", x"25",
	x"27", x"26", x"24", x"24", x"22", x"20", x"21", x"1D", x"19", x"19", x"0D", x"0A",
	x"07", x"03", x"F9", x"FA", x"F4", x"F2", x"F0", x"EA", x"EC", x"EC", x"E9", x"E7",
	x"E6", x"E6", x"E5", x"E8", x"E7", x"E5", x"E7", x"E1", x"E5", x"E7", x"E7", x"E6",
	x"E5", x"EC", x"EB", x"ED", x"EF", x"F4", x"F8", x"FF", x"04", x"06", x"0E", x"0E",
	x"15", x"17", x"1E", x"20", x"24", x"27", x"26", x"26", x"21", x"26", x"20", x"21",
	x"1F", x"1F", x"1C", x"19", x"19", x"0F", x"0F", x"06", x"FA", x"F6", x"ED", x"E7",
	x"E1", x"E1", x"DA", x"DB", x"DA", x"D6", x"D5", x"D6", x"D7", x"DB", x"E2", x"E2",
	x"E5", x"E9", x"EC", x"F1", x"F3", x"FA", x"02", x"01", x"05", x"04", x"04", x"08",
	x"07", x"0F", x"0F", x"13", x"0D", x"0C", x"0A", x"0D", x"13", x"16", x"14", x"1B",
	x"1A", x"16", x"16", x"16", x"18", x"18", x"1A", x"1C", x"18", x"15", x"11", x"0C",
	x"07", x"01", x"00", x"FB", x"F6", x"F2", x"EA", x"E6", x"E2", x"E0", x"DE", x"DA",
	x"D8", x"D6", x"DB", x"DC", x"DB", x"D8", x"DE", x"DF", x"E2", x"E7", x"EB", x"F4",
	x"F8", x"01", x"06", x"0C", x"0F", x"14", x"13", x"17", x"1C", x"1D", x"20", x"20",
	x"1D", x"22", x"1F", x"1F", x"1E", x"18", x"17", x"13", x"10", x"0B", x"0A", x"05",
	x"00", x"FE", x"FE", x"FE", x"FB", x"F8", x"F9", x"FA", x"FA", x"FB", x"F9", x"F6",
	x"F5", x"F3", x"F0", x"EE", x"EA", x"EA", x"E4", x"E4", x"E0", x"DD", x"E0", x"DE",
	x"DF", x"E1", x"E5", x"E8", x"EE", x"F2", x"FB", x"FC", x"01", x"05", x"0A", x"0F",
	x"10", x"12", x"18", x"1A", x"1C", x"1D", x"23", x"23", x"25", x"26", x"23", x"22",
	x"1E", x"1B", x"14", x"14", x"0B", x"04", x"03", x"FE", x"FA", x"F7", x"F4", x"F3",
	x"F0", x"EF", x"EB", x"E9", x"EA", x"E6", x"EA", x"E6", x"E6", x"E9", x"E7", x"E9",
	x"E8", x"EA", x"E9", x"ED", x"F4", x"F3", x"F7", x"F9", x"F9", x"FD", x"FA", x"FF",
	x"FD", x"FF", x"02", x"01", x"03", x"07", x"08", x"0C", x"10", x"11", x"12", x"16",
	x"19", x"1A", x"1B", x"21", x"1E", x"1D", x"1E", x"1C", x"19", x"15", x"10", x"0A",
	x"04", x"00", x"F9", x"F5", x"F4", x"F0", x"EC", x"EF", x"E8", x"E9", x"E3", x"E2",
	x"E2", x"E1", x"E5", x"E7", x"E9", x"EE", x"EF", x"EE", x"EE", x"EF", x"F0", x"F4",
	x"F7", x"FA", x"FE", x"FF", x"01", x"02", x"04", x"07", x"08", x"08", x"0A", x"0E",
	x"10", x"12", x"15", x"12", x"14", x"14", x"12", x"17", x"15", x"14", x"14", x"11",
	x"0F", x"0C", x"0B", x"0C", x"0C", x"0A", x"08", x"06", x"02", x"FC", x"F9", x"F7",
	x"F2", x"F2", x"E9", x"E8", x"E4", x"E2", x"E2", x"E1", x"E0", x"E2", x"E5", x"E7",
	x"EA", x"EB", x"EE", x"F0", x"F4", x"F6", x"FB", x"FC", x"FC", x"01", x"04", x"06",
	x"0A", x"0F", x"13", x"13", x"15", x"16", x"15", x"16", x"11", x"12", x"11", x"0F",
	x"0E", x"10", x"10", x"0F", x"0C", x"0B", x"0B", x"06", x"04", x"04", x"01", x"03",
	x"04", x"00", x"02", x"FF", x"FD", x"F8", x"F6", x"F3", x"EF", x"ED", x"E7", x"E7",
	x"E6", x"E5", x"E7", x"E6", x"E9", x"EC", x"EC", x"EE", x"ED", x"EF", x"EF", x"F0",
	x"F1", x"F5", x"FA", x"FD", x"04", x"07", x"0C", x"10", x"0F", x"15", x"16", x"1A",
	x"1B", x"1B", x"1B", x"19", x"1A", x"19", x"18", x"15", x"14", x"0E", x"0B", x"08",
	x"04", x"00", x"FB", x"F8", x"F6", x"F5", x"F5", x"F6", x"F6", x"F7", x"F3", x"F5",
	x"F6", x"F2", x"F3", x"F1", x"EF", x"F3", x"F2", x"F1", x"F1", x"EE", x"F0", x"EC",
	x"EE", x"EF", x"EF", x"F2", x"F1", x"F4", x"F4", x"F6", x"F8", x"FA", x"01", x"03",
	x"07", x"0D", x"10", x"13", x"12", x"13", x"14", x"15", x"16", x"17", x"19", x"1A",
	x"19", x"1B", x"19", x"15", x"15", x"0E", x"0B", x"04", x"00", x"F9", x"F4", x"F1",
	x"F0", x"F0", x"F0", x"F0", x"F1", x"F0", x"F1", x"EC", x"ED", x"EB", x"EC", x"EB",
	x"ED", x"ED", x"EF", x"F0", x"F2", x"F3", x"F4", x"F5", x"F8", x"FA", x"F9", x"FE",
	x"FE", x"01", x"03", x"04", x"07", x"08", x"08", x"0A", x"09", x"0D", x"0D", x"0B",
	x"0C", x"0C", x"0C", x"0C", x"10", x"11", x"11", x"12", x"14", x"16", x"15", x"12",
	x"0F", x"0B", x"07", x"03", x"01", x"FF", x"FB", x"F9", x"F5", x"F3", x"EC", x"EB",
	x"E9", x"E7", x"E5", x"E4", x"E2", x"E3", x"E5", x"E8", x"EB", x"ED", x"F0", x"F2",
	x"F6", x"F7", x"FD", x"00", x"02", x"05", x"07", x"09", x"08", x"0B", x"0C", x"0B",
	x"0D", x"0E", x"0D", x"0E", x"0D", x"0D", x"0B", x"0A", x"08", x"07", x"06", x"08",
	x"08", x"0B", x"0C", x"0C", x"0C", x"0C", x"0D", x"08", x"06", x"04", x"02", x"FE",
	x"FE", x"FC", x"F9", x"F9", x"F5", x"F4", x"F0", x"EE", x"ED", x"E9", x"E8", x"E7",
	x"E8", x"E8", x"EA", x"EC", x"EC", x"ED", x"EF", x"F0", x"F5", x"F6", x"F8", x"FD",
	x"FD", x"02", x"06", x"0A", x"0D", x"12", x"15", x"15", x"19", x"18", x"1A", x"17",
	x"18", x"16", x"14", x"13", x"0E", x"0C", x"07", x"04", x"FE", x"FF", x"FC", x"FB",
	x"FC", x"FA", x"FB", x"F8", x"F9", x"F8", x"F7", x"F6", x"F9", x"F7", x"F8", x"F8",
	x"F8", x"F9", x"F6", x"F5", x"F4", x"F4", x"F2", x"F1", x"F1", x"F0", x"F0", x"F2",
	x"EF", x"F2", x"F3", x"F6", x"F8", x"F6", x"FA", x"FB", x"FE", x"04", x"04", x"0A",
	x"0C", x"0D", x"11", x"13", x"14", x"15", x"18", x"17", x"18", x"16", x"15", x"16",
	x"12", x"10", x"0E", x"0A", x"08", x"03", x"FF", x"FA", x"F8", x"F4", x"F3", x"EF",
	x"EF", x"EE", x"ED", x"ED", x"EC", x"EF", x"EE", x"EF", x"EE", x"EF", x"EF", x"F0",
	x"F3", x"F4", x"F7", x"FA", x"FB", x"FE", x"FF", x"01", x"01", x"01", x"00", x"01",
	x"01", x"02", x"02", x"02", x"02", x"05", x"05", x"07", x"06", x"08", x"09", x"0A",
	x"0C", x"0F", x"10", x"11", x"10", x"11", x"11", x"11", x"0F", x"0E", x"0A", x"08",
	x"04", x"02", x"FE", x"FC", x"F8", x"F7", x"F6", x"F2", x"F2", x"F0", x"EE", x"ED",
	x"EB", x"EB", x"EB", x"EC", x"EB", x"EE", x"EC", x"EF", x"F0", x"F3", x"F4", x"F8",
	x"FB", x"00", x"02", x"03", x"05", x"06", x"07", x"09", x"0B", x"0A", x"0B", x"0C",
	x"0D", x"0B", x"0D", x"0C", x"0C", x"0B", x"0B", x"0A", x"0B", x"0A", x"09", x"08",
	x"07", x"08", x"05", x"03", x"03", x"01", x"02", x"00", x"FE", x"FE", x"FB", x"FC",
	x"F9", x"F8", x"F6", x"F4", x"F3", x"F2", x"F1", x"EF", x"EF", x"ED", x"EE", x"EE",
	x"EE", x"F0", x"F2", x"F3", x"F4", x"F7", x"FA", x"FA", x"FE", x"FE", x"01", x"04",
	x"06", x"09", x"0C", x"0C", x"0F", x"10", x"0F", x"10", x"0E", x"0E", x"0E", x"0E",
	x"0B", x"0B", x"08", x"07", x"04", x"05", x"02", x"05", x"03", x"02", x"03", x"00",
	x"00", x"FD", x"FD", x"FC", x"FD", x"FB", x"FB", x"F9", x"FA", x"F7", x"F5", x"F3",
	x"F3", x"F1", x"F0", x"EF", x"F1", x"F0", x"F1", x"F0", x"F1", x"F2", x"F3", x"F5",
	x"F6", x"F9", x"F9", x"FD", x"00", x"04", x"06", x"08", x"0B", x"0D", x"0E", x"0F",
	x"11", x"13", x"11", x"11", x"0F", x"0F", x"0D", x"0D", x"0A", x"0A", x"07", x"07",
	x"02", x"01", x"FF", x"FF", x"FB", x"FB", x"F9", x"F9", x"F7", x"F8", x"F6", x"F6",
	x"F6", x"F5", x"F6", x"F5", x"F7", x"F7", x"F7", x"F9", x"FB", x"F9", x"FB", x"F9",
	x"FA", x"F8", x"F9", x"F8", x"F9", x"F9", x"F8", x"FA", x"F8", x"F8", x"FA", x"F9",
	x"FD", x"FF", x"01", x"03", x"06", x"07", x"0B", x"0C", x"0D", x"0F", x"0E", x"11",
	x"11", x"13", x"13", x"11", x"12", x"11", x"0E", x"0B", x"08", x"03", x"FF", x"FB",
	x"F9", x"F6", x"F4", x"F2", x"F0", x"EE", x"EF", x"ED", x"EF", x"EE", x"F1", x"F1",
	x"F3", x"F4", x"F6", x"F6", x"F8", x"F9", x"FA", x"FD", x"FC", x"FE", x"FF", x"01",
	x"01", x"02", x"03", x"05", x"05", x"06", x"05", x"05", x"04", x"04", x"03", x"03",
	x"02", x"02", x"02", x"03", x"04", x"03", x"04", x"04", x"07", x"08", x"09", x"09",
	x"0C", x"0A", x"0B", x"09", x"08", x"07", x"04", x"04", x"01", x"01", x"FE", x"FB",
	x"FA", x"F6", x"F4", x"F0", x"F0", x"ED", x"EC", x"EB", x"EB", x"EA", x"EB", x"EB",
	x"EE", x"F0", x"F3", x"F7", x"FA", x"FF", x"02", x"06", x"07", x"09", x"0A", x"0C",
	x"0B", x"0D", x"0C", x"0D", x"0D", x"0C", x"0B", x"09", x"08", x"06", x"05", x"04",
	x"04", x"04", x"04", x"04", x"02", x"02", x"00", x"01", x"FF", x"FE", x"FE", x"FD",
	x"FC", x"FC", x"FB", x"FC", x"FC", x"FD", x"FC", x"FE", x"FE", x"FC", x"FC", x"FA",
	x"F7", x"F7", x"F6", x"F4", x"F4", x"F3", x"F4", x"F4", x"F5", x"F4", x"F7", x"F6",
	x"F8", x"F7", x"FA", x"FB", x"FC", x"FF", x"00", x"04", x"05", x"09", x"0B", x"0D",
	x"0F", x"10", x"12", x"12", x"12", x"11", x"0F", x"0D", x"0B", x"09", x"06", x"04",
	x"01", x"01", x"FD", x"FC", x"FA", x"F8", x"F6", x"F7", x"F5", x"F6", x"F5", x"F7",
	x"F6", x"F7", x"F8", x"F6", x"F7", x"F6", x"F8", x"F7", x"F7", x"FA", x"F9", x"FB",
	x"FB", x"FB", x"FD", x"FD", x"FC", x"FC", x"FD", x"FB", x"FD", x"FE", x"FF", x"FF",
	x"01", x"02", x"03", x"05", x"06", x"08", x"09", x"0B", x"0B", x"0A", x"0C", x"0B",
	x"0A", x"0A", x"09", x"0A", x"07", x"07", x"07", x"05", x"04", x"01", x"01", x"FE",
	x"FD", x"FB", x"F9", x"F8", x"F7", x"F6", x"F5", x"F4", x"F5", x"F4", x"F4", x"F4",
	x"F3", x"F4", x"F4", x"F4", x"F6", x"F7", x"F9", x"FA", x"FD", x"FC", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"01", x"01", x"02", x"02", x"04", x"04", x"07", x"06", x"08",
	x"08", x"09", x"09", x"08", x"09", x"08", x"09", x"08", x"09", x"07", x"08", x"07",
	x"07", x"05", x"05", x"03", x"01", x"FF", x"FE", x"FB", x"F8", x"F8", x"F6", x"F5",
	x"F5", x"F4", x"F2", x"F4", x"F2", x"F3", x"F3", x"F4", x"F4", x"F6", x"F6", x"F8",
	x"F8", x"FA", x"FA", x"FE", x"FF", x"00", x"03", x"04", x"04", x"05", x"04", x"06",
	x"06", x"06", x"05", x"05", x"04", x"05", x"04", x"05", x"05", x"05", x"05", x"06",
	x"05", x"06", x"05", x"05", x"06", x"05", x"06", x"05", x"05", x"04", x"02", x"02",
	x"FF", x"FD", x"FE", x"FB", x"FB", x"FA", x"F8", x"F8", x"F5", x"F5", x"F3", x"F3",
	x"F1", x"F2", x"F1", x"F0", x"F1", x"F0", x"F3", x"F4", x"F6", x"F7", x"FB", x"FC",
	x"00", x"01", x"04", x"06", x"09", x"0A", x"0D", x"0C", x"0E", x"0E", x"0E", x"0D",
	x"0D", x"0A", x"0A", x"07", x"06", x"04", x"03", x"01", x"00", x"FE", x"FE", x"FC",
	x"FD", x"FB", x"FC", x"FC", x"FB", x"FC", x"FC", x"FD", x"FD", x"FC", x"FE", x"FC",
	x"FE", x"FD", x"FD", x"FE", x"FC", x"FC", x"FB", x"F9", x"F8", x"F6", x"F5", x"F6",
	x"F4", x"F5", x"F6", x"F4", x"F7", x"F7", x"F9", x"FB", x"FB", x"FE", x"FE", x"02",
	x"02", x"05", x"07", x"0A", x"0A", x"0D", x"0D", x"0F", x"0F", x"10", x"11", x"0F",
	x"0F", x"0C", x"0B", x"09", x"07", x"04", x"03", x"FF", x"FC", x"FB", x"F7", x"F6",
	x"F4", x"F2", x"F2", x"F1", x"F1", x"F1", x"F2", x"F4", x"F3", x"F5", x"F7", x"F9",
	x"FB", x"FB", x"FD", x"FE", x"00", x"01", x"02", x"03", x"03", x"03", x"03", x"01",
	x"01", x"FF", x"FF", x"FE", x"FF", x"FD", x"FE", x"FE", x"00", x"FF", x"01", x"01",
	x"02", x"04", x"04", x"08", x"08", x"0A", x"0A", x"0A", x"0B", x"09", x"0A", x"08",
	x"09", x"07", x"06", x"04", x"02", x"FF", x"FE", x"FB", x"FA", x"F8", x"F6", x"F3",
	x"F3", x"F2", x"F1", x"F1", x"F0", x"F1", x"F1", x"F3", x"F4", x"F4", x"F6", x"F7",
	x"FA", x"FB", x"FF", x"01", x"02", x"04", x"05", x"07", x"07", x"09", x"08", x"0A",
	x"09", x"09", x"08", x"08", x"06", x"07", x"05", x"05", x"03", x"03", x"01", x"02",
	x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"00", x"FE", x"FE", x"FC", x"FD", x"FC", x"FA", x"FA", x"F8", x"F7", x"F6",
	x"F4", x"F5", x"F3", x"F4", x"F5", x"F5", x"F7", x"F6", x"F9", x"F9", x"FC", x"FF",
	x"FF", x"03", x"04", x"05", x"07", x"07", x"09", x"0A", x"09", x"0B", x"0A", x"0A",
	x"0A", x"09", x"07", x"07", x"04", x"05", x"03", x"03", x"01", x"02", x"00", x"01",
	x"FE", x"FF", x"FD", x"FC", x"FB", x"FB", x"F9", x"FA", x"F9", x"FA", x"FA", x"F9",
	x"FB", x"F9", x"FA", x"F9", x"FA", x"F9", x"F9", x"F8", x"F8", x"F8", x"F7", x"F9",
	x"F9", x"FB", x"FC", x"FD", x"FD", x"00", x"00", x"01", x"01", x"03", x"04", x"04",
	x"06", x"07", x"06", x"08", x"07", x"09", x"09", x"0A", x"08", x"09", x"08", x"06",
	x"05", x"03", x"03", x"01", x"00", x"FE", x"FE", x"FC", x"FB", x"FB", x"F9", x"FA",
	x"F9", x"F8", x"FA", x"F9", x"FA", x"F9", x"FA", x"F9", x"FB", x"FB", x"FB", x"FC",
	x"FB", x"FC", x"FC", x"FD", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD",
	x"FD", x"FD", x"FE", x"FD", x"FF", x"00", x"02", x"03", x"05", x"05", x"07", x"08",
	x"0A", x"0A", x"0B", x"0B", x"09", x"09", x"07", x"07", x"06", x"04", x"04", x"01",
	x"00", x"FF", x"FC", x"FB", x"F9", x"F8", x"F7", x"F6", x"F6", x"F5", x"F5", x"F4",
	x"F6", x"F5", x"F6", x"F8", x"F8", x"F9", x"F9", x"FC", x"FC", x"FF", x"00", x"01",
	x"02", x"03", x"04", x"04", x"03", x"04", x"03", x"04", x"02", x"02", x"00", x"01",
	x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"01", x"01", x"01", x"02", x"03",
	x"02", x"04", x"03", x"05", x"04", x"06", x"05", x"05", x"06", x"04", x"04", x"02",
	x"FF", x"FE", x"FA", x"FA", x"F8", x"F5", x"F5", x"F4", x"F3", x"F3", x"F2", x"F4",
	x"F3", x"F4", x"F5", x"F7", x"F7", x"FA", x"FC", x"FD", x"01", x"01", x"04", x"05",
	x"07", x"08", x"0A", x"09", x"0A", x"09", x"09", x"08", x"06", x"07", x"04", x"04",
	x"04", x"03", x"01", x"00", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FE", x"FE", x"FC", x"FC", x"F9", x"F9", x"F7", x"F7", x"F7",
	x"F6", x"F7", x"F8", x"F9", x"FB", x"FB", x"FE", x"FF", x"02", x"03", x"05", x"05",
	x"08", x"08", x"09", x"0A", x"0A", x"0B", x"0A", x"0B", x"09", x"09", x"06", x"06",
	x"03", x"02", x"00", x"FE", x"FD", x"FB", x"FA", x"FA", x"F8", x"F8", x"F7", x"F8",
	x"F7", x"F8", x"F9", x"F8", x"FA", x"FB", x"FB", x"FD", x"FE", x"FE", x"FF", x"FE",
	x"FF", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"01", x"01", x"00", x"02", x"01", x"03", x"03",
	x"05", x"04", x"06", x"05", x"07", x"06", x"07", x"05", x"06", x"05", x"03", x"03",
	x"01", x"01", x"FE", x"FE", x"FC", x"FB", x"FA", x"F7", x"F7", x"F6", x"F7", x"F6",
	x"F7", x"F7", x"F7", x"F8", x"F8", x"FA", x"FB", x"FB", x"FD", x"FD", x"FF", x"FF",
	x"01", x"01", x"02", x"03", x"02", x"03", x"02", x"03", x"02", x"01", x"02", x"01",
	x"01", x"00", x"01", x"02", x"01", x"03", x"02", x"04", x"04", x"04", x"03", x"05",
	x"03", x"04", x"02", x"02", x"01", x"01", x"00", x"00", x"FE", x"FF", x"FF", x"FD",
	x"FD", x"FB", x"FC", x"FA", x"FA", x"F8", x"F8", x"F8", x"F7", x"F8", x"F7", x"F9",
	x"FA", x"FA", x"FA", x"FC", x"FC", x"FE", x"FF", x"FF", x"01", x"01", x"02", x"03",
	x"03", x"04", x"03", x"04", x"04", x"03", x"04", x"03", x"04", x"02", x"03", x"02",
	x"03", x"03", x"01", x"02", x"02", x"00", x"01", x"FF", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FD", x"FD", x"FC",
	x"FB", x"FA", x"F9", x"F9", x"F8", x"F8", x"F7", x"F8", x"F8", x"F8", x"FA", x"FA",
	x"FC", x"FC", x"FE", x"FE", x"00", x"00", x"02", x"02", x"05", x"06", x"05", x"07",
	x"07", x"08", x"08", x"07", x"08", x"06", x"06", x"04", x"03", x"02", x"00", x"00",
	x"FE", x"FE", x"FC", x"FD", x"FB", x"FC", x"FB", x"FC", x"FB", x"FC", x"FC", x"FD",
	x"FC", x"FD", x"FD", x"FE", x"FE", x"FD", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FC", x"FD", x"FB", x"FC", x"FA", x"FB", x"FA", x"FB", x"FA", x"FC", x"FD",
	x"FD", x"FE", x"FF", x"FF", x"01", x"02", x"04", x"04", x"06", x"07", x"06", x"08",
	x"07", x"08", x"08", x"06", x"07", x"06", x"06", x"04", x"03", x"02", x"00", x"FF",
	x"FD", x"FC", x"FB", x"F9", x"F8", x"F6", x"F7", x"F5", x"F7", x"F6", x"F8", x"F7",
	x"FA", x"FA", x"FB", x"FC", x"FE", x"FE", x"00", x"00", x"02", x"02", x"02", x"03",
	x"02", x"02", x"02", x"00", x"01", x"FF", x"00", x"FF", x"00", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"00", x"01", x"00", x"02", x"02", x"03", x"04", x"04", x"05",
	x"05", x"06", x"05", x"06", x"04", x"04", x"02", x"02", x"01", x"FE", x"FE", x"FD",
	x"FC", x"FB", x"F9", x"F9", x"F8", x"F7", x"F7", x"F6", x"F7", x"F6", x"F8", x"F8",
	x"F8", x"FA", x"FB", x"FC", x"FE", x"FE", x"00", x"02", x"02", x"04", x"04", x"05",
	x"06", x"05", x"06", x"06", x"04", x"05", x"04", x"03", x"03", x"01", x"02", x"02",
	x"00", x"00", x"FE", x"FF", x"FF", x"FD", x"FE", x"FD", x"FF", x"FE", x"00", x"FF",
	x"01", x"00", x"01", x"01", x"00", x"01", x"FF", x"00", x"FE", x"FE", x"FD", x"FD",
	x"FB", x"FB", x"F9", x"F9", x"F9", x"F8", x"F9", x"F9", x"F8", x"F9", x"F9", x"FB",
	x"FC", x"FC", x"FE", x"FF", x"01", x"01", x"03", x"03", x"05", x"04", x"06", x"05",
	x"06", x"06", x"06", x"05", x"06", x"05", x"05", x"03", x"03", x"01", x"01", x"FF",
	x"FF", x"FD", x"FD", x"FC", x"FD", x"FC", x"FC", x"FB", x"FC", x"FD", x"FC", x"FD",
	x"FC", x"FD", x"FC", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FD", x"FE", x"FD",
	x"FD", x"FC", x"FC", x"FC", x"FB", x"FC", x"FB", x"FC", x"FB", x"FD", x"FE", x"FE",
	x"00", x"FF", x"01", x"01", x"03", x"02", x"04", x"04", x"06", x"06", x"07", x"06",
	x"07", x"06", x"06", x"05", x"05", x"03", x"03", x"01", x"FF", x"FE", x"FD", x"FB",
	x"FB", x"FA", x"FA", x"FA", x"F9", x"F9", x"F9", x"FA", x"FA", x"FB", x"FA", x"FC",
	x"FC", x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FE",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"02", x"02", x"04", x"03", x"05", x"04", x"06", x"05", x"05",
	x"04", x"04", x"03", x"02", x"02", x"00", x"00", x"FE", x"FD", x"FD", x"FB", x"FB",
	x"F9", x"F9", x"F8", x"F8", x"F7", x"F8", x"F7", x"F9", x"F8", x"FA", x"FA", x"FC",
	x"FC", x"FE", x"FF", x"FF", x"01", x"01", x"03", x"03", x"04", x"05", x"04", x"05",
	x"04", x"04", x"03", x"03", x"02", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FE", x"00", x"FF", x"01", x"01", x"00", x"01", x"00", x"02", x"01", x"02", x"02",
	x"01", x"02", x"01", x"02", x"00", x"01", x"00", x"FD", x"FD", x"FB", x"FA", x"F8",
	x"F9", x"F7", x"F8", x"F7", x"F8", x"F8", x"F9", x"F9", x"FB", x"FB", x"FD", x"FD",
	x"FF", x"00", x"00", x"02", x"03", x"03", x"05", x"05", x"05", x"06", x"06", x"05",
	x"05", x"04", x"04", x"03", x"03", x"02", x"02", x"01", x"00", x"00", x"FE", x"FE",
	x"FD", x"FD", x"FB", x"FC", x"FB", x"FC", x"FB", x"FD", x"FC", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FD",
	x"FC", x"FC", x"FB", x"FC", x"FB", x"FB", x"FB", x"FB", x"FC", x"FC", x"FE", x"FF",
	x"FF", x"01", x"01", x"03", x"03", x"05", x"04", x"06", x"06", x"07", x"07", x"07",
	x"06", x"05", x"05", x"04", x"02", x"01", x"00", x"FD", x"FD", x"FC", x"FA", x"FB",
	x"FA", x"FB", x"FA", x"FB", x"FB", x"FC", x"FB", x"FC", x"FC", x"FC", x"FD", x"FC",
	x"FE", x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"01",
	x"00", x"02", x"02", x"02", x"03", x"02", x"04", x"03", x"04", x"03", x"04", x"04",
	x"03", x"03", x"01", x"02", x"00", x"00", x"FE", x"FD", x"FC", x"FA", x"FB", x"FA",
	x"FA", x"F8", x"F9", x"F8", x"F9", x"F9", x"FA", x"FA", x"FC", x"FC", x"FE", x"FE",
	x"00", x"01", x"01", x"02", x"02", x"02", x"02", x"02", x"02", x"01", x"02", x"01",
	x"01", x"01", x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"02", x"01", x"02", x"01", x"02", x"02", x"00",
	x"01", x"FF", x"FF", x"FF", x"FD", x"FD", x"FC", x"FC", x"FC", x"FA", x"FB", x"F9",
	x"FA", x"F9", x"FA", x"FA", x"FA", x"FA", x"FB", x"FB", x"FD", x"FD", x"FF", x"FF",
	x"01", x"01", x"03", x"03", x"04", x"04", x"05", x"06", x"05", x"05", x"04", x"04",
	x"04", x"02", x"02", x"01", x"FF", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FC", x"FD", x"FC", x"FA", x"FB",
	x"FB", x"FA", x"FB", x"FA", x"FC", x"FC", x"FC", x"FE", x"FE", x"00", x"01", x"00",
	x"02", x"03", x"02", x"04", x"04", x"05", x"05", x"06", x"06", x"05", x"04", x"05",
	x"03", x"03", x"02", x"02", x"00", x"FF", x"FE", x"FC", x"FC", x"FB", x"FA", x"FA",
	x"F9", x"FA", x"FB", x"FA", x"FB", x"FB", x"FD", x"FC", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"FE", x"FF", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FF", x"FF", x"00",
	x"00", x"02", x"02", x"03", x"03", x"04", x"05", x"04", x"05", x"04", x"04", x"03",
	x"03", x"01", x"01", x"FF", x"FE", x"FE", x"FC", x"FC", x"FB", x"FB", x"FA", x"FA",
	x"F9", x"FA", x"F9", x"FA", x"F9", x"FB", x"FB", x"FB", x"FD", x"FD", x"FE", x"FE",
	x"00", x"01", x"01", x"02", x"03", x"02", x"03", x"02", x"03", x"02", x"01", x"02",
	x"00", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"FF",
	x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"01",
	x"00", x"00", x"00", x"FE", x"FE", x"FD", x"FD", x"FB", x"FC", x"FA", x"FB", x"FA",
	x"FB", x"FA", x"FB", x"FA", x"FC", x"FC", x"FC", x"FD", x"FD", x"FF", x"FE", x"00",
	x"01", x"01", x"03", x"02", x"04", x"04", x"03", x"04", x"03", x"04", x"03", x"02",
	x"02", x"00", x"01", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FD", x"FE", x"FE", x"FF", x"FE", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FE", x"FF", x"FD", x"FE", x"FC", x"FD", x"FB", x"FC", x"FC", x"FB", x"FC",
	x"FB", x"FC", x"FC", x"FD", x"FE", x"FD", x"FF", x"FF", x"00", x"00", x"02", x"02",
	x"03", x"03", x"04", x"04", x"04", x"04", x"03", x"04", x"02", x"03", x"02", x"01",
	x"01", x"FF", x"FF", x"FF", x"FD", x"FE", x"FD", x"FC", x"FD", x"FB", x"FC", x"FB",
	x"FD", x"FD", x"FC", x"FE", x"FD", x"FE", x"FE", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FC", x"FD",
	x"FC", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"00", x"01", x"00", x"02", x"02",
	x"03", x"04", x"04", x"05", x"05", x"04", x"05", x"04", x"04", x"02", x"02", x"00",
	x"00", x"FF", x"FE", x"FC", x"FC", x"FA", x"FB", x"FA", x"FA", x"FA", x"FA", x"FA",
	x"FB", x"FC", x"FC", x"FD", x"FC", x"FE", x"FE", x"00", x"FF", x"01", x"00", x"02",
	x"01", x"02", x"01", x"02", x"01", x"01", x"00", x"01", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"02", x"03", x"02", x"04", x"03", x"04", x"02", x"03", x"03", x"02", x"01", x"00",
	x"00", x"FE", x"FE", x"FE", x"FC", x"FC", x"FB", x"FA", x"FA", x"F9", x"F9", x"F8",
	x"FA", x"F9", x"FB", x"FB", x"FB", x"FD", x"FE", x"FF", x"01", x"01", x"03", x"03",
	x"04", x"04", x"05", x"04", x"04", x"03", x"04", x"02", x"03", x"02", x"01", x"00",
	x"00", x"FF", x"FD", x"FE", x"FC", x"FD", x"FC", x"FD", x"FE", x"FE", x"FE", x"FF",
	x"FE", x"00", x"FF", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FD", x"FD", x"FB", x"FC", x"FC", x"FA", x"FB", x"FA",
	x"FC", x"FB", x"FC", x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"02", x"03",
	x"03", x"04", x"04", x"04", x"04", x"04", x"03", x"04", x"02", x"03", x"01", x"01",
	x"FF", x"00", x"FF", x"FE", x"FE", x"FD", x"FD", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FC", x"FD", x"FC", x"FE", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"01",
	x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"02", x"01", x"03",
	x"03", x"03", x"02", x"03", x"02", x"03", x"03", x"01", x"02", x"00", x"01", x"00",
	x"FE", x"FF", x"FD", x"FD", x"FC", x"FC", x"FC", x"FB", x"FC", x"FB", x"FD", x"FD",
	x"FC", x"FE", x"FD", x"FE", x"FD", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"01", x"01", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FE",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"01", x"00", x"01", x"01", x"02",
	x"01", x"03", x"02", x"03", x"01", x"02", x"01", x"01", x"FF", x"00", x"FE", x"FE",
	x"FC", x"FD", x"FC", x"FC", x"FB", x"FC", x"FC", x"FB", x"FC", x"FB", x"FC", x"FC",
	x"FC", x"FD", x"FD", x"FF", x"FE", x"00", x"00", x"01", x"01", x"02", x"02", x"03",
	x"02", x"02", x"01", x"02", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"01", x"00",
	x"01", x"00", x"01", x"01", x"00", x"01", x"01", x"FF", x"00", x"FF", x"FF", x"FE",
	x"FE", x"FD", x"FC", x"FC", x"FB", x"FB", x"FA", x"FB", x"FB", x"FB", x"FC", x"FB",
	x"FD", x"FD", x"FE", x"FF", x"FF", x"01", x"02", x"01", x"03", x"04", x"04", x"03",
	x"04", x"03", x"04", x"03", x"03", x"02", x"02", x"01", x"FF", x"00", x"FE", x"FE",
	x"FE", x"FC", x"FD", x"FB", x"FC", x"FD", x"FC", x"FD", x"FD", x"FE", x"FE", x"FF",
	x"00", x"FF", x"00", x"00", x"01", x"00", x"01", x"01", x"00", x"00", x"FF", x"00",
	x"FF", x"FE", x"FE", x"FD", x"FD", x"FD", x"FC", x"FD", x"FB", x"FD", x"FC", x"FD",
	x"FC", x"FE", x"FD", x"FF", x"FF", x"00", x"01", x"02", x"02", x"03", x"03", x"04",
	x"03", x"04", x"04", x"03", x"04", x"02", x"03", x"01", x"01", x"FF", x"FF", x"FE",
	x"FE", x"FC", x"FC", x"FB", x"FB", x"FA", x"FB", x"FB", x"FA", x"FB", x"FC", x"FB",
	x"FD", x"FD", x"FE", x"FE", x"00", x"00", x"01", x"01", x"02", x"01", x"02", x"01",
	x"01", x"00", x"01", x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FE", x"FD", x"FE",
	x"FD", x"FD", x"FF", x"FE", x"FF", x"FE", x"00", x"00", x"01", x"00", x"02", x"01",
	x"02", x"02", x"03", x"03", x"02", x"02", x"01", x"01", x"00", x"00", x"FE", x"FF",
	x"FD", x"FD", x"FD", x"FB", x"FC", x"FB", x"FB", x"FA", x"FB", x"FB", x"FC", x"FB",
	x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"02", x"02", x"02",
	x"03", x"02", x"03", x"02", x"02", x"01", x"01", x"00", x"00", x"00", x"FE", x"FF",
	x"FD", x"FE", x"FD", x"FE", x"FD", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE",
	x"FF", x"FD", x"FE", x"FC", x"FD", x"FC", x"FD", x"FC", x"FD", x"FC", x"FD", x"FC",
	x"FE", x"FD", x"FF", x"FE", x"00", x"01", x"00", x"02", x"01", x"03", x"03", x"03",
	x"02", x"03", x"02", x"02", x"01", x"01", x"00", x"00", x"FF", x"00", x"FE", x"FF",
	x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FE", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FC", x"FD", x"FC", x"FD", x"FC", x"FE", x"FD", x"FE", x"FE", x"FF",
	x"00", x"FF", x"01", x"00", x"01", x"01", x"02", x"01", x"02", x"01", x"03", x"03",
	x"02", x"02", x"01", x"02", x"00", x"01", x"FF", x"00", x"FF", x"FE", x"FE", x"FC",
	x"FD", x"FD", x"FC", x"FC", x"FD", x"FC", x"FD", x"FD", x"FD", x"FE", x"FF", x"FE",
	x"FF", x"00", x"FF", x"00", x"00", x"01", x"00", x"01", x"00", x"00", x"00", x"FF",
	x"00", x"FE", x"FF", x"FF", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FF",
	x"FE", x"00", x"FF", x"01", x"01", x"01", x"02", x"02", x"03", x"02", x"03", x"02",
	x"03", x"01", x"02", x"01", x"01", x"00", x"FF", x"FF", x"FD", x"FD", x"FC", x"FC",
	x"FB", x"FB", x"FA", x"FB", x"FA", x"FC", x"FB", x"FD", x"FC", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"01", x"00", x"01", x"01", x"02", x"01", x"02", x"02", x"01", x"02",
	x"01", x"00", x"01", x"FF", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FD", x"FE", x"FD", x"FF", x"FE", x"00", x"00", x"00", x"01", x"02", x"01", x"02",
	x"01", x"02", x"01", x"02", x"00", x"01", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD",
	x"FB", x"FC", x"FB", x"FB", x"FA", x"FA", x"FC", x"FB", x"FC", x"FC", x"FD", x"FE",
	x"FF", x"00", x"01", x"01", x"02", x"03", x"02", x"04", x"03", x"04", x"04", x"02",
	x"03", x"01", x"01", x"01", x"FF", x"00", x"FE", x"FF", x"FE", x"FE", x"FD", x"FD",
	x"FC", x"FD", x"FC", x"FD", x"FD", x"FE", x"FD", x"FF", x"FF", x"FE", x"00", x"00",
	x"FF", x"01", x"00", x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"FF", x"FE",
	x"FE", x"FD", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD", x"FC", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"02", x"02", x"02", x"03", x"03", x"03", x"03", x"03",
	x"03", x"03", x"02", x"02", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD",
	x"FD", x"FC", x"FC", x"FC", x"FD", x"FD", x"FC", x"FE", x"FD", x"FD", x"FF", x"FE",
	x"00", x"FF", x"01", x"00", x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"FE",
	x"FF", x"FF", x"FE", x"FF", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"00", x"FF", x"01", x"01", x"01", x"01", x"02", x"02", x"02", x"02", x"01",
	x"02", x"00", x"01", x"FF", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FC", x"FD",
	x"FD", x"FC", x"FD", x"FC", x"FD", x"FC", x"FD", x"FD", x"FE", x"FE", x"FF", x"00",
	x"FF", x"00", x"00", x"01", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01",
	x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FC", x"FD",
	x"FB", x"FD", x"FC", x"FD", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"00", x"FF",
	x"01", x"01", x"00", x"02", x"02", x"01", x"02", x"01", x"02", x"01", x"01", x"01",
	x"00", x"00", x"00", x"FE", x"FF", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD",
	x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"01", x"00",
	x"01", x"00", x"00", x"FF", x"FF", x"00", x"FE", x"FF", x"FE", x"FD", x"FD", x"FC",
	x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FD", x"FE", x"FF", x"FE", x"00", x"01",
	x"01", x"01", x"02", x"02", x"03", x"02", x"03", x"02", x"03", x"01", x"02", x"00",
	x"01", x"FF", x"00", x"FE", x"FF", x"FD", x"FE", x"FC", x"FD", x"FD", x"FC", x"FD",
	x"FC", x"FD", x"FD", x"FD", x"FE", x"FD", x"FF", x"FF", x"FF", x"00", x"01", x"01",
	x"00", x"01", x"00", x"01", x"01", x"00", x"00", x"00", x"FE", x"FF", x"FD", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE", x"FF", x"FE", x"00",
	x"FF", x"01", x"00", x"01", x"01", x"02", x"01", x"03", x"02", x"03", x"02", x"01",
	x"02", x"00", x"01", x"00", x"FF", x"FE", x"FE", x"FD", x"FD", x"FB", x"FC", x"FB",
	x"FC", x"FB", x"FC", x"FD", x"FC", x"FE", x"FD", x"FF", x"FF", x"FF", x"00", x"FF",
	x"01", x"00", x"02", x"02", x"01", x"02", x"01", x"01", x"00", x"01", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FF", x"FE", x"FF",
	x"FE", x"00", x"FF", x"00", x"00", x"01", x"01", x"00", x"02", x"00", x"01", x"00",
	x"01", x"01", x"FF", x"00", x"FE", x"FF", x"FD", x"FE", x"FD", x"FD", x"FC", x"FD",
	x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FD", x"FE", x"FE", x"FF", x"00", x"00",
	x"01", x"00", x"02", x"01", x"02", x"01", x"02", x"02", x"02", x"00", x"01", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FD", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FE", x"FD", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"01", x"00", x"02", x"01", x"02", x"02", x"01", x"02", x"02", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FE", x"FE", x"FF", x"FE", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"FF", x"01", x"00",
	x"01", x"01", x"02", x"01", x"02", x"02", x"01", x"02", x"00", x"01", x"01", x"FF",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FC", x"FD", x"FC", x"FC", x"FD",
	x"FC", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"00", x"01", x"01",
	x"01", x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FE",
	x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FE", x"FE", x"FF", x"FE", x"00", x"FF",
	x"01", x"01", x"01", x"02", x"01", x"02", x"01", x"02", x"00", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"FE", x"FD", x"FD", x"FC", x"FD", x"FC", x"FB", x"FC", x"FD",
	x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"FE", x"00", x"FF", x"01", x"01", x"00",
	x"02", x"02", x"02", x"01", x"02", x"01", x"02", x"01", x"01", x"01", x"FF", x"FF",
	x"FE", x"FE", x"FD", x"FE", x"FE", x"FC", x"FE", x"FD", x"FE", x"FD", x"FF", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01",
	x"00", x"00", x"FF", x"FF", x"FE", x"FD", x"FE", x"FD", x"FC", x"FD", x"FC", x"FD",
	x"FD", x"FC", x"FD", x"FD", x"FE", x"FF", x"FE", x"00", x"FF", x"01", x"00", x"02",
	x"01", x"02", x"02", x"01", x"02", x"01", x"02", x"01", x"01", x"01", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FD", x"FE", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"01", x"00", x"01", x"00",
	x"01", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FE", x"FE", x"FD", x"FF", x"FE", x"00", x"00", x"FF", x"01", x"00",
	x"02", x"01", x"02", x"02", x"01", x"02", x"02", x"00", x"01", x"00", x"00", x"00",
	x"FE", x"FF", x"FD", x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FD", x"FC", x"FE",
	x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"01", x"00", x"01", x"00",
	x"01", x"00", x"01", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"01", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FD", x"FE", x"FC", x"FD", x"FC", x"FC", x"FD", x"FC", x"FE",
	x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"FF", x"01", x"01", x"00", x"01", x"00",
	x"01", x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FE",
	x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"FF", x"FE", x"FF", x"00", x"FF", x"00",
	x"00", x"01", x"00", x"01", x"00", x"01", x"01", x"FF", x"00", x"FF", x"00", x"FE",
	x"FF", x"FD", x"FE", x"FD", x"FE", x"FE", x"FC", x"FD", x"FC", x"FD", x"FD", x"FE",
	x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"00", x"01", x"01", x"02", x"01",
	x"02", x"01", x"02", x"01", x"01", x"00", x"01", x"FF", x"00", x"FE", x"FF", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"00", x"FF", x"01", x"00", x"01", x"00", x"01", x"01", x"00", x"00", x"FF",
	x"00", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FE", x"FF", x"FE", x"00", x"FF", x"01", x"01", x"00", x"02", x"01",
	x"02", x"01", x"02", x"01", x"02", x"00", x"01", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FD", x"FE", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FF", x"FE", x"00", x"FF", x"01", x"00", x"01", x"01", x"00", x"01", x"01",
	x"00", x"01", x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FD", x"FE", x"FE", x"FF", x"FF", x"FE", x"00", x"00", x"FF", x"01", x"00", x"01",
	x"01", x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"FF", x"00", x"FF", x"FF",
	x"FE", x"FE", x"FD", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"01", x"01", x"01", x"00", x"01", x"00",
	x"01", x"01", x"00", x"01", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF",
	x"FD", x"FE", x"FE", x"FD", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"FF", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"01", x"00", x"01", x"00", x"02", x"01",
	x"02", x"00", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FD", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FD", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FF",
	x"FE", x"FF", x"00", x"FF", x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"01",
	x"00", x"01", x"00", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"00",
	x"00", x"FF", x"00", x"01", x"01", x"01", x"00", x"01", x"01", x"00", x"00", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FD", x"FE", x"FD", x"FD", x"FE", x"FD", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"01", x"01", x"00", x"01", x"00",
	x"02", x"00", x"01", x"00", x"01", x"00", x"FF", x"FF", x"FE", x"FF", x"FD", x"FE",
	x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FD", x"FD", x"FE", x"FD", x"FE", x"FF",
	x"FE", x"00", x"00", x"00", x"01", x"00", x"02", x"01", x"02", x"00", x"01", x"00",
	x"01", x"00", x"FF", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FD", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"01", x"00", x"01",
	x"00", x"01", x"01", x"00", x"01", x"01", x"00", x"00", x"00", x"FE", x"FF", x"FD",
	x"FE", x"FE", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FE", x"FD", x"FE", x"FE",
	x"FF", x"FF", x"00", x"FF", x"01", x"01", x"00", x"02", x"01", x"02", x"02", x"01",
	x"01", x"00", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD",
	x"FC", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"FF", x"01",
	x"00", x"01", x"01", x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"FE", x"FF",
	x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE", x"FD", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"01", x"01", x"00", x"01", x"01", x"02", x"02",
	x"00", x"01", x"00", x"01", x"00", x"00", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FF", x"FF", x"FE", x"00",
	x"FF", x"00", x"01", x"00", x"01", x"00", x"01", x"01", x"00", x"00", x"00", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"00", x"FF", x"00", x"00", x"01", x"01", x"00", x"01", x"00", x"01",
	x"00", x"01", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"00", x"00",
	x"FF", x"00", x"00", x"FF", x"01", x"01", x"00", x"01", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"01", x"01", x"00", x"01",
	x"01", x"00", x"00", x"FF", x"FF", x"00", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"00", x"FF",
	x"00", x"01", x"01", x"01", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"FF",
	x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD",
	x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"01", x"00", x"01",
	x"00", x"01", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"FD", x"FE",
	x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"00",
	x"FF", x"01", x"01", x"01", x"00", x"02", x"01", x"02", x"01", x"01", x"01", x"01",
	x"00", x"FF", x"00", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"01", x"00",
	x"01", x"00", x"01", x"00", x"01", x"FF", x"00", x"FF", x"00", x"FE", x"FE", x"FF",
	x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"FE",
	x"00", x"00", x"FF", x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"01",
	x"00", x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FD", x"FE", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF",
	x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"01", x"00", x"01", x"00", x"01", x"00",
	x"01", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"00",
	x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00",
	x"00", x"FF", x"FE", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"00",
	x"FF", x"01", x"00", x"01", x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FD", x"FE", x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"01", x"01",
	x"01", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"00",
	x"FF", x"00", x"FF", x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"FF",
	x"00", x"00", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"01",
	x"01", x"00", x"01", x"00", x"01", x"01", x"00", x"00", x"FF", x"00", x"FF", x"FE",
	x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"01",
	x"00", x"01", x"00", x"02", x"01", x"00", x"01", x"00", x"01", x"FF", x"00", x"FF",
	x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"01", x"01", x"00", x"01",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FD", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"01", x"00", x"01", x"01", x"01", x"00", x"01", x"00", x"00", x"FF",
	x"00", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"00", x"01",
	x"00", x"00", x"01", x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FD", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"00", x"00", x"00",
	x"00", x"00", x"01", x"01", x"01", x"00", x"01", x"FF", x"00", x"00", x"FF", x"00",
	x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"01", x"00", x"01",
	x"01", x"01", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FE",
	x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"01", x"00", x"01", x"00", x"01", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE", x"FD", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"01", x"00", x"01", x"01",
	x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"01", x"00", x"01", x"00", x"01", x"FF", x"00",
	x"00", x"00", x"00", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FD", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"00",
	x"01", x"00", x"01", x"00", x"01", x"01", x"FF", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"FF", x"00", x"01", x"00", x"01", x"00", x"01", x"01", x"01",
	x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE",
	x"FF", x"FE", x"00", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"01",
	x"00", x"01", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"01", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FF", x"FE",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"01", x"01", x"00",
	x"01", x"00", x"01", x"FF", x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FE", x"FF", x"FE", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"01", x"00",
	x"01", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FD", x"FE", x"FD", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"01", x"01", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF",
	x"00", x"FF", x"00", x"00", x"FF", x"01", x"00", x"01", x"01", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FD", x"FE", x"FD",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FF",
	x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF",
	x"FE", x"00", x"00", x"FF", x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"00",
	x"01", x"FF", x"FF", x"00", x"FF", x"00", x"FE", x"FE", x"FF", x"FE", x"FE", x"FD",
	x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00",
	x"FF", x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"00", x"01", x"00", x"01",
	x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"00",
	x"01", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"FE", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"00",
	x"FF", x"00", x"00", x"FF", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"00",
	x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"00", x"FF", x"00", x"00", x"00", x"01",
	x"01", x"01", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF", x"FE", x"00",
	x"FF", x"00", x"00", x"FF", x"01", x"01", x"00", x"01", x"00", x"01", x"00", x"00",
	x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"FF",
	x"01", x"00", x"00", x"01", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"01", x"00", x"01", x"01", x"00", x"01", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FD", x"FE",
	x"FE", x"FD", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"01", x"00", x"00", x"01", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"01", x"01", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FE", x"FF", x"FE", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"01", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FD", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"01",
	x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FE",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FD", x"FD", x"FE", x"FD", x"FF", x"FE",
	x"FF", x"FE", x"FE", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"FF",
	x"01", x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"01", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FD", x"FF", x"FE", x"FF", x"FE", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FD", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FF", x"FE", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"01", x"01",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE"
	);
	
signal cnt_out: unsigned(14 downto 0) := (others => '0');	
signal play_sound: std_logic := '0';
constant cnt_max: integer := 8959;
signal out_signal: signed(7 downto 0) := x"00";

begin
	
process (CLK)
begin
    if rising_edge(CLK) then
        if RST = '1' then
            play_sound <= '0';
        elsif PLAY = '1' then
            play_sound <= '1';
        elsif PLAY = '0' and cnt_out = cnt_max then
            play_sound <= '0';
        end if;
    end if;
end process;

	
-- 12bit counter
process (CLK)
begin     
    if rising_edge(CLK) then
        if RST = '1' then
            cnt_out <= (others => '0');
        elsif CE = '1' and play_sound = '1' then
            cnt_out <= cnt_out + 1;       
        end if;
        if cnt_out = cnt_max then
            cnt_out <= (others => '0');            
        end if;        
    end if;
end process;

process (CLK) 
begin
    if rising_edge(CLK) then
        if RST = '1' then
            out_signal <= x"00";
        elsif CE = '1' then
            out_signal <= tom1_sound(conv_integer(cnt_out));
        end if;
    end if;    
end process;

SAMPLE_OUT <= out_signal;

end Behavioral;