----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 25.12.2018 17:39:59
-- Design Name: 
-- Module Name: HHat - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity HHat is
    Port ( CLK : in STD_LOGIC;
           CE : in STD_LOGIC;
           RST : in STD_LOGIC;
           PLAY : in STD_LOGIC;
           SAMPLE_OUT : out signed(7 downto 0)
           );
end HHat;

architecture Behavioral of HHat is

type memory is array (0 to 8857) of signed(7 downto 0);
constant hhat_sound: memory := (
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"01", x"00", x"01", x"02", x"01", x"00", x"02", x"03",
	x"FC", x"03", x"FD", x"E7", x"FF", x"02", x"EB", x"C7", x"AE", x"CE", x"CD", x"D7",
	x"E5", x"EA", x"1C", x"40", x"32", x"0A", x"FB", x"14", x"2E", x"F7", x"DE", x"EA",
	x"18", x"2D", x"FF", x"EA", x"FD", x"3C", x"2C", x"03", x"EB", x"0D", x"1C", x"E7",
	x"EB", x"11", x"14", x"02", x"E9", x"CF", x"E8", x"18", x"08", x"26", x"28", x"24",
	x"2C", x"03", x"1F", x"25", x"F1", x"08", x"2F", x"35", x"10", x"D7", x"D4", x"F3",
	x"07", x"24", x"FB", x"D6", x"F1", x"F6", x"EE", x"EC", x"0E", x"12", x"10", x"1C",
	x"FE", x"DB", x"E3", x"09", x"1E", x"20", x"1C", x"08", x"20", x"F7", x"DD", x"07",
	x"EA", x"CF", x"C1", x"E5", x"F4", x"DA", x"CD", x"D4", x"B8", x"E8", x"0C", x"DD",
	x"EA", x"0A", x"F0", x"CD", x"D0", x"EA", x"DF", x"E7", x"1C", x"21", x"EE", x"BD",
	x"D9", x"1F", x"0A", x"09", x"0F", x"E6", x"E1", x"F0", x"F4", x"CF", x"D9", x"DC",
	x"D9", x"ED", x"0D", x"07", x"B3", x"D7", x"18", x"0C", x"00", x"16", x"11", x"D7",
	x"EF", x"22", x"0D", x"F7", x"FB", x"F5", x"CA", x"D4", x"E2", x"BC", x"CA", x"E6",
	x"E4", x"D0", x"CE", x"EB", x"E3", x"E2", x"05", x"1D", x"17", x"E7", x"C7", x"DE",
	x"EA", x"E3", x"D1", x"C5", x"DC", x"07", x"00", x"D2", x"DA", x"FE", x"03", x"04",
	x"2A", x"1A", x"E2", x"16", x"2B", x"2E", x"35", x"06", x"E5", x"01", x"08", x"F0",
	x"06", x"E6", x"E1", x"EA", x"0D", x"00", x"E6", x"D4", x"E6", x"EF", x"F2", x"F4",
	x"DF", x"D4", x"FA", x"23", x"27", x"00", x"F1", x"05", x"FA", x"03", x"09", x"E7",
	x"F0", x"2B", x"16", x"10", x"29", x"24", x"18", x"12", x"2E", x"1A", x"1D", x"2B",
	x"25", x"21", x"EC", x"E7", x"D7", x"CF", x"DB", x"CA", x"AA", x"D7", x"24", x"E7",
	x"D2", x"E0", x"A2", x"BC", x"DC", x"E9", x"FA", x"F4", x"FB", x"08", x"F0", x"ED",
	x"1B", x"23", x"0D", x"ED", x"0E", x"21", x"01", x"01", x"14", x"13", x"1F", x"FA",
	x"D9", x"09", x"28", x"E7", x"DA", x"0A", x"16", x"18", x"F9", x"F5", x"28", x"07",
	x"F3", x"E9", x"09", x"36", x"30", x"08", x"ED", x"08", x"09", x"08", x"28", x"03",
	x"0D", x"06", x"F5", x"0E", x"DE", x"06", x"01", x"EB", x"E8", x"F9", x"1F", x"06",
	x"CA", x"C8", x"DD", x"C1", x"AE", x"EB", x"FD", x"C8", x"9A", x"CD", x"E7", x"C0",
	x"BB", x"9D", x"BE", x"01", x"F6", x"18", x"06", x"F1", x"2C", x"03", x"ED", x"1E",
	x"23", x"39", x"2E", x"2F", x"0C", x"E7", x"FC", x"3C", x"1B", x"1B", x"1C", x"06",
	x"2C", x"1A", x"08", x"F2", x"EB", x"0A", x"17", x"36", x"2B", x"22", x"1E", x"17",
	x"1E", x"E1", x"DE", x"17", x"18", x"D8", x"E7", x"EB", x"FB", x"36", x"22", x"07",
	x"22", x"32", x"02", x"E9", x"16", x"2A", x"2E", x"13", x"23", x"43", x"32", x"18",
	x"17", x"11", x"32", x"41", x"38", x"2C", x"04", x"FF", x"23", x"2B", x"21", x"14",
	x"17", x"27", x"0C", x"EA", x"E7", x"EA", x"12", x"06", x"CF", x"D1", x"FC", x"F8",
	x"EB", x"05", x"E6", x"D1", x"D1", x"07", x"34", x"F8", x"E3", x"F6", x"E6", x"EC",
	x"05", x"02", x"F1", x"FC", x"EB", x"EE", x"D5", x"CB", x"DF", x"F8", x"26", x"EA",
	x"B5", x"F3", x"FC", x"F9", x"11", x"27", x"09", x"CF", x"E3", x"43", x"0E", x"DF",
	x"F8", x"00", x"E4", x"C9", x"CE", x"CE", x"E8", x"22", x"0E", x"1C", x"33", x"2C",
	x"F1", x"E4", x"FA", x"15", x"15", x"04", x"2C", x"12", x"DF", x"F6", x"13", x"39",
	x"22", x"29", x"15", x"F0", x"02", x"E3", x"0F", x"4C", x"21", x"12", x"0C", x"2A",
	x"25", x"E4", x"D0", x"EC", x"0A", x"FC", x"D5", x"02", x"35", x"23", x"1A", x"24",
	x"2F", x"33", x"25", x"04", x"16", x"3D", x"21", x"FE", x"12", x"1C", x"34", x"21",
	x"CD", x"D5", x"E5", x"FB", x"09", x"FE", x"44", x"30", x"1E", x"31", x"17", x"2D",
	x"2C", x"2C", x"58", x"3D", x"0F", x"C9", x"B6", x"F7", x"1F", x"0F", x"13", x"F4",
	x"0B", x"31", x"17", x"E5", x"EA", x"1C", x"27", x"2E", x"2D", x"30", x"FF", x"09",
	x"2B", x"11", x"30", x"2D", x"1C", x"20", x"28", x"05", x"D4", x"0C", x"2D", x"1C",
	x"F1", x"0A", x"FD", x"E1", x"D8", x"0B", x"3B", x"08", x"D4", x"14", x"FD", x"20",
	x"F6", x"B8", x"0A", x"0B", x"1F", x"0B", x"16", x"FD", x"02", x"08", x"F4", x"F1",
	x"27", x"16", x"E6", x"E4", x"E8", x"F8", x"F4", x"F4", x"CF", x"F8", x"F7", x"03",
	x"F8", x"F8", x"27", x"13", x"1F", x"3C", x"04", x"DF", x"F3", x"0B", x"04", x"DF",
	x"BE", x"01", x"39", x"1D", x"FA", x"D9", x"DD", x"F5", x"FF", x"0C", x"29", x"13",
	x"DE", x"D2", x"F9", x"3B", x"47", x"35", x"F5", x"F1", x"2A", x"DB", x"11", x"16",
	x"EC", x"31", x"40", x"1E", x"17", x"19", x"03", x"F2", x"F8", x"23", x"1C", x"31",
	x"0C", x"22", x"25", x"28", x"28", x"0F", x"1A", x"2B", x"2D", x"24", x"31", x"0D",
	x"EF", x"25", x"33", x"0D", x"1E", x"3C", x"38", x"3E", x"09", x"09", x"03", x"F7",
	x"F9", x"05", x"18", x"1E", x"33", x"25", x"19", x"06", x"EB", x"E8", x"02", x"0C",
	x"FD", x"C2", x"D4", x"13", x"1E", x"FD", x"FB", x"E6", x"CF", x"E6", x"16", x"18",
	x"F2", x"FC", x"04", x"FD", x"FC", x"F9", x"F9", x"16", x"EF", x"00", x"1F", x"F6",
	x"00", x"EF", x"E3", x"E6", x"DB", x"DF", x"EB", x"01", x"EF", x"EC", x"EA", x"FE",
	x"10", x"07", x"1D", x"09", x"BF", x"D2", x"15", x"20", x"22", x"E2", x"FB", x"24",
	x"26", x"19", x"0F", x"06", x"E2", x"0B", x"30", x"22", x"04", x"F9", x"04", x"13",
	x"15", x"09", x"0C", x"25", x"E9", x"E6", x"E4", x"1A", x"33", x"FF", x"FB", x"F6",
	x"06", x"EB", x"C5", x"2C", x"3B", x"29", x"22", x"0B", x"04", x"1B", x"30", x"09",
	x"F4", x"1A", x"13", x"F3", x"0B", x"26", x"28", x"27", x"34", x"04", x"D7", x"19",
	x"16", x"EC", x"DA", x"FF", x"EA", x"09", x"01", x"F3", x"DF", x"E6", x"ED", x"C5",
	x"E8", x"08", x"F4", x"18", x"02", x"FA", x"CB", x"E3", x"1C", x"06", x"10", x"F1",
	x"E4", x"D1", x"FD", x"0E", x"ED", x"25", x"1D", x"FF", x"D7", x"DC", x"FA", x"10",
	x"1B", x"12", x"28", x"0B", x"E4", x"F5", x"F1", x"DF", x"DD", x"11", x"39", x"FA",
	x"F7", x"D6", x"DD", x"EB", x"CC", x"08", x"31", x"38", x"07", x"B9", x"E3", x"F3",
	x"FC", x"1D", x"30", x"0C", x"E1", x"E6", x"C4", x"DF", x"FD", x"E1", x"02", x"06",
	x"F2", x"D6", x"F3", x"1D", x"FD", x"E4", x"E9", x"D1", x"E4", x"E7", x"FA", x"D9",
	x"BC", x"DD", x"D1", x"E0", x"0B", x"2A", x"27", x"21", x"E9", x"B2", x"DA", x"13",
	x"FD", x"F1", x"EF", x"E8", x"E6", x"03", x"09", x"1D", x"39", x"12", x"04", x"01",
	x"F8", x"29", x"1D", x"02", x"E4", x"16", x"29", x"1B", x"F5", x"F0", x"34", x"41",
	x"36", x"1F", x"12", x"1A", x"0E", x"0D", x"01", x"02", x"E8", x"FB", x"24", x"0F",
	x"EA", x"E0", x"09", x"17", x"1E", x"2A", x"1F", x"05", x"F6", x"F0", x"17", x"1A",
	x"15", x"15", x"0C", x"D1", x"EA", x"EE", x"13", x"2E", x"12", x"18", x"27", x"10",
	x"E7", x"E6", x"1C", x"1E", x"E8", x"14", x"0A", x"03", x"F4", x"EF", x"2D", x"0F",
	x"0F", x"2F", x"28", x"07", x"D9", x"B2", x"C5", x"E6", x"1B", x"1C", x"FA", x"0C",
	x"14", x"EB", x"D4", x"07", x"F6", x"0A", x"0C", x"09", x"02", x"02", x"EA", x"DD",
	x"EE", x"F9", x"1B", x"34", x"14", x"EE", x"D4", x"02", x"F6", x"EF", x"03", x"EB",
	x"FE", x"0B", x"D9", x"F4", x"FE", x"06", x"EE", x"FC", x"32", x"28", x"E3", x"D7",
	x"C1", x"D9", x"0C", x"16", x"1D", x"06", x"EC", x"F4", x"FB", x"C1", x"C3", x"29",
	x"0F", x"BB", x"E3", x"24", x"31", x"02", x"D2", x"E5", x"EC", x"16", x"11", x"15",
	x"16", x"09", x"F1", x"FB", x"17", x"E6", x"DF", x"FE", x"08", x"1A", x"24", x"06",
	x"1D", x"DC", x"D2", x"10", x"05", x"2A", x"16", x"E3", x"D7", x"C8", x"E4", x"0D",
	x"0A", x"19", x"0B", x"F6", x"E3", x"08", x"EB", x"0B", x"3D", x"10", x"F3", x"EF",
	x"F0", x"D3", x"A1", x"BC", x"0E", x"29", x"17", x"06", x"D9", x"D2", x"E6", x"09",
	x"1B", x"37", x"0E", x"D8", x"03", x"1C", x"E8", x"FD", x"08", x"0C", x"20", x"26",
	x"DF", x"AA", x"FB", x"0F", x"16", x"12", x"FB", x"EB", x"DC", x"01", x"F6", x"EC",
	x"FC", x"07", x"17", x"2A", x"0D", x"CE", x"E3", x"0D", x"00", x"E5", x"FE", x"F0",
	x"E1", x"FB", x"0C", x"0E", x"F3", x"CB", x"EC", x"0B", x"00", x"DF", x"CD", x"ED",
	x"00", x"1D", x"2F", x"0A", x"11", x"04", x"EC", x"E5", x"EF", x"E9", x"0C", x"1F",
	x"1D", x"27", x"F6", x"EF", x"D6", x"E2", x"00", x"27", x"13", x"FD", x"0C", x"18",
	x"01", x"FB", x"23", x"17", x"2E", x"33", x"FF", x"DF", x"C7", x"D9", x"0A", x"29",
	x"16", x"F8", x"04", x"18", x"09", x"04", x"01", x"FE", x"F8", x"0C", x"FD", x"B9",
	x"BD", x"E5", x"E3", x"0B", x"1E", x"FC", x"E7", x"F4", x"10", x"EE", x"DB", x"E5",
	x"E2", x"EA", x"E7", x"E1", x"E0", x"D6", x"FA", x"12", x"17", x"EB", x"EE", x"DF",
	x"B7", x"FF", x"FB", x"DF", x"E5", x"EC", x"0E", x"C1", x"E2", x"0D", x"F6", x"F0",
	x"F6", x"02", x"0F", x"05", x"D5", x"D5", x"E4", x"08", x"01", x"D6", x"0F", x"EF",
	x"F2", x"1B", x"00", x"F1", x"E6", x"BA", x"DD", x"F6", x"FD", x"08", x"E3", x"F0",
	x"14", x"05", x"2B", x"F1", x"C0", x"D7", x"16", x"F8", x"C5", x"0F", x"33", x"ED",
	x"CF", x"E3", x"FA", x"FD", x"1A", x"20", x"01", x"0B", x"03", x"EF", x"DC", x"EC",
	x"E7", x"D8", x"F5", x"FA", x"0B", x"24", x"08", x"C7", x"D3", x"06", x"FC", x"FB",
	x"F8", x"F7", x"D6", x"E6", x"10", x"07", x"E4", x"E2", x"CF", x"FF", x"0A", x"F7",
	x"E6", x"DA", x"05", x"FF", x"E8", x"E5", x"FC", x"24", x"27", x"0F", x"E8", x"F0",
	x"01", x"1A", x"07", x"FD", x"1D", x"19", x"EB", x"B6", x"02", x"1D", x"EA", x"EA",
	x"F5", x"18", x"11", x"E7", x"D7", x"FF", x"0D", x"04", x"E6", x"E7", x"1E", x"26",
	x"F5", x"E0", x"F7", x"EB", x"0A", x"1D", x"F8", x"C7", x"AB", x"ED", x"01", x"08",
	x"17", x"F1", x"FE", x"D4", x"C4", x"DC", x"EB", x"F3", x"F8", x"E7", x"E9", x"F9",
	x"1C", x"EA", x"B6", x"DD", x"2D", x"1D", x"DE", x"DB", x"07", x"09", x"CB", x"E1",
	x"DF", x"08", x"06", x"CE", x"EE", x"0A", x"14", x"EA", x"E1", x"FD", x"01", x"F4",
	x"F1", x"08", x"F2", x"E1", x"01", x"14", x"FB", x"FA", x"08", x"D8", x"FA", x"2F",
	x"0B", x"D9", x"D8", x"08", x"3B", x"F4", x"D6", x"F0", x"DB", x"FC", x"18", x"19",
	x"11", x"F7", x"DF", x"DC", x"F8", x"EA", x"07", x"EE", x"DD", x"15", x"26", x"11",
	x"EB", x"01", x"0E", x"E2", x"CB", x"03", x"29", x"19", x"E2", x"EB", x"08", x"D8",
	x"DA", x"F3", x"14", x"04", x"D6", x"CC", x"E7", x"FA", x"31", x"F4", x"D3", x"0F",
	x"1B", x"09", x"E4", x"DC", x"F9", x"F0", x"19", x"13", x"E1", x"D4", x"21", x"25",
	x"CA", x"D8", x"F6", x"F0", x"CC", x"E5", x"02", x"DF", x"E4", x"F4", x"F7", x"02",
	x"D5", x"C9", x"C4", x"11", x"2F", x"13", x"04", x"F3", x"EE", x"ED", x"D4", x"FD",
	x"0A", x"12", x"10", x"FA", x"11", x"1A", x"F5", x"0A", x"17", x"E3", x"E3", x"29",
	x"21", x"18", x"1F", x"33", x"05", x"07", x"0E", x"F7", x"E9", x"E5", x"16", x"16",
	x"10", x"15", x"22", x"28", x"F7", x"F5", x"11", x"0D", x"24", x"20", x"04", x"0F",
	x"25", x"28", x"07", x"EC", x"F5", x"23", x"26", x"01", x"D4", x"11", x"13", x"E5",
	x"10", x"07", x"EB", x"10", x"1B", x"06", x"DF", x"D8", x"04", x"F4", x"0B", x"12",
	x"F9", x"0A", x"FC", x"C9", x"DB", x"FB", x"FA", x"F2", x"0D", x"EF", x"C6", x"B4",
	x"E2", x"FE", x"0E", x"F0", x"D9", x"0C", x"03", x"E9", x"F2", x"BB", x"E2", x"FB",
	x"D8", x"EA", x"FD", x"14", x"FF", x"CE", x"DD", x"F7", x"03", x"F9", x"CF", x"DF",
	x"E1", x"06", x"2E", x"04", x"D7", x"C9", x"F2", x"FB", x"01", x"E1", x"FB", x"02",
	x"E8", x"0F", x"26", x"00", x"EC", x"12", x"08", x"0C", x"F3", x"E4", x"FA", x"F0",
	x"10", x"15", x"0D", x"12", x"01", x"F2", x"EB", x"08", x"23", x"1C", x"23", x"04",
	x"EC", x"D9", x"CF", x"2D", x"13", x"F4", x"EF", x"0A", x"12", x"05", x"10", x"EF",
	x"FD", x"27", x"05", x"F7", x"16", x"17", x"DE", x"D9", x"11", x"35", x"35", x"F8",
	x"CA", x"E3", x"06", x"FF", x"FF", x"13", x"FD", x"12", x"02", x"09", x"15", x"17",
	x"0B", x"F3", x"F5", x"1D", x"33", x"17", x"FD", x"FA", x"FB", x"16", x"FE", x"E2",
	x"FE", x"03", x"16", x"03", x"DB", x"EE", x"22", x"22", x"21", x"1F", x"0A", x"FF",
	x"05", x"1A", x"22", x"FE", x"DC", x"E8", x"1D", x"FC", x"FB", x"1A", x"2A", x"00",
	x"F3", x"04", x"02", x"F4", x"E8", x"13", x"2B", x"22", x"0B", x"EE", x"07", x"10",
	x"07", x"0F", x"E5", x"CE", x"DB", x"28", x"1B", x"11", x"18", x"1D", x"08", x"FA",
	x"0D", x"F7", x"F4", x"E0", x"E7", x"0B", x"12", x"19", x"11", x"1A", x"F2", x"CF",
	x"F4", x"02", x"F2", x"FF", x"0E", x"0D", x"E5", x"DF", x"08", x"D5", x"E7", x"05",
	x"F0", x"DE", x"FD", x"11", x"03", x"E1", x"EB", x"13", x"06", x"05", x"F6", x"04",
	x"F9", x"C4", x"F4", x"11", x"15", x"05", x"EA", x"D1", x"D6", x"CD", x"DF", x"14",
	x"13", x"F9", x"FD", x"15", x"1B", x"E6", x"DA", x"F7", x"FC", x"F1", x"04", x"FD",
	x"ED", x"D0", x"E7", x"08", x"11", x"EC", x"E8", x"1D", x"1B", x"ED", x"DC", x"E3",
	x"CF", x"FB", x"33", x"FC", x"EC", x"DD", x"F5", x"F2", x"E8", x"01", x"1A", x"F9",
	x"FC", x"06", x"E2", x"EA", x"04", x"0D", x"EE", x"10", x"23", x"07", x"D6", x"00",
	x"F9", x"F4", x"FC", x"08", x"28", x"0D", x"ED", x"E9", x"06", x"0E", x"18", x"14",
	x"02", x"13", x"1A", x"18", x"12", x"17", x"03", x"EF", x"EF", x"09", x"19", x"19",
	x"13", x"07", x"22", x"13", x"14", x"18", x"FE", x"00", x"01", x"1F", x"2C", x"F9",
	x"E8", x"F1", x"14", x"10", x"0F", x"E5", x"DB", x"0F", x"04", x"06", x"15", x"1E",
	x"0C", x"FA", x"1C", x"0E", x"F7", x"EE", x"0C", x"05", x"03", x"0E", x"12", x"0E",
	x"01", x"F1", x"FF", x"E9", x"E9", x"F4", x"08", x"17", x"F5", x"02", x"16", x"13",
	x"0A", x"E2", x"03", x"0B", x"0F", x"F9", x"E0", x"04", x"0A", x"08", x"02", x"08",
	x"0D", x"00", x"02", x"F8", x"01", x"27", x"1D", x"1E", x"0F", x"09", x"07", x"06",
	x"11", x"00", x"F9", x"16", x"20", x"19", x"10", x"E9", x"CC", x"FC", x"24", x"15",
	x"09", x"0E", x"FD", x"E3", x"DF", x"0D", x"30", x"17", x"F4", x"F2", x"FA", x"12",
	x"FB", x"FD", x"F7", x"F5", x"FA", x"F1", x"FE", x"E7", x"DF", x"03", x"0B", x"12",
	x"14", x"06", x"01", x"FC", x"E2", x"EB", x"DF", x"DE", x"FF", x"07", x"16", x"FA",
	x"F1", x"F4", x"F9", x"F0", x"F5", x"F0", x"12", x"0B", x"03", x"07", x"0B", x"03",
	x"FA", x"03", x"0F", x"04", x"EA", x"D7", x"F7", x"0A", x"02", x"F5", x"FA", x"03",
	x"E3", x"E8", x"FD", x"0C", x"1A", x"0D", x"19", x"08", x"E7", x"D2", x"D1", x"FA",
	x"11", x"01", x"07", x"FC", x"E2", x"F5", x"E6", x"E9", x"0C", x"0A", x"FC", x"EB",
	x"FA", x"EE", x"E4", x"EE", x"0C", x"0D", x"03", x"06", x"F5", x"FC", x"0E", x"06",
	x"F2", x"F8", x"01", x"15", x"0E", x"08", x"FF", x"FC", x"16", x"17", x"07", x"F3",
	x"05", x"29", x"1A", x"0D", x"1B", x"2B", x"15", x"01", x"FF", x"19", x"25", x"1B",
	x"1F", x"25", x"12", x"05", x"07", x"13", x"17", x"F1", x"0C", x"23", x"0E", x"FA",
	x"0A", x"18", x"09", x"F6", x"13", x"1D", x"12", x"32", x"1E", x"0C", x"05", x"04",
	x"01", x"06", x"0F", x"09", x"FE", x"0A", x"04", x"F4", x"E5", x"EA", x"E6", x"F3",
	x"1B", x"10", x"FC", x"F3", x"08", x"13", x"08", x"DD", x"D2", x"05", x"14", x"FE",
	x"F5", x"FF", x"08", x"01", x"F7", x"F7", x"F7", x"09", x"F1", x"EF", x"F3", x"13",
	x"1A", x"F5", x"03", x"06", x"FB", x"F8", x"11", x"0F", x"E4", x"D9", x"EF", x"0C",
	x"01", x"0D", x"05", x"02", x"FD", x"F5", x"F2", x"E7", x"E4", x"F9", x"0F", x"0D",
	x"E2", x"F7", x"04", x"F3", x"FD", x"FE", x"1A", x"F2", x"F8", x"17", x"0F", x"04",
	x"F6", x"FC", x"02", x"01", x"F5", x"F2", x"10", x"12", x"13", x"1B", x"0F", x"F9",
	x"F9", x"04", x"F9", x"F3", x"16", x"19", x"FD", x"01", x"05", x"F4", x"F0", x"04",
	x"0A", x"FF", x"F9", x"06", x"09", x"EA", x"FE", x"FA", x"FE", x"12", x"04", x"EB",
	x"FB", x"13", x"0C", x"F3", x"06", x"14", x"0B", x"17", x"17", x"FE", x"0A", x"00",
	x"F2", x"F3", x"F8", x"06", x"03", x"0C", x"0F", x"0A", x"10", x"0A", x"FE", x"01",
	x"1E", x"08", x"0C", x"0D", x"F0", x"FB", x"00", x"03", x"03", x"11", x"1C", x"0C",
	x"0C", x"FB", x"F4", x"06", x"03", x"0E", x"07", x"EF", x"EF", x"F7", x"17", x"13",
	x"04", x"0E", x"F8", x"05", x"F9", x"0B", x"16", x"14", x"20", x"14", x"06", x"E9",
	x"E9", x"06", x"0B", x"1E", x"04", x"07", x"13", x"FB", x"03", x"08", x"FD", x"15",
	x"07", x"1A", x"FE", x"EC", x"14", x"11", x"03", x"01", x"F9", x"0C", x"02", x"F3",
	x"FD", x"F9", x"11", x"02", x"FE", x"10", x"07", x"EE", x"EB", x"07", x"04", x"06",
	x"0E", x"F2", x"F4", x"F5", x"FA", x"E7", x"E2", x"04", x"02", x"F2", x"F5", x"02",
	x"0B", x"F8", x"FB", x"F2", x"F3", x"01", x"FD", x"FD", x"0A", x"F6", x"E8", x"F2",
	x"04", x"FA", x"EF", x"E6", x"EE", x"13", x"12", x"FB", x"FB", x"00", x"03", x"0B",
	x"09", x"FF", x"07", x"FF", x"01", x"0B", x"04", x"01", x"03", x"04", x"0C", x"12",
	x"FE", x"FA", x"F9", x"0C", x"15", x"22", x"10", x"F8", x"FD", x"FF", x"10", x"1D",
	x"0F", x"04", x"F7", x"12", x"01", x"0D", x"17", x"07", x"0C", x"05", x"0A", x"0C",
	x"02", x"0C", x"14", x"14", x"02", x"EC", x"EB", x"F8", x"08", x"10", x"FC", x"F5",
	x"F6", x"0B", x"13", x"03", x"F7", x"F6", x"F7", x"FB", x"FA", x"FD", x"F5", x"FC",
	x"08", x"03", x"FD", x"E8", x"DD", x"F3", x"FF", x"0A", x"00", x"FC", x"09", x"EE",
	x"ED", x"01", x"02", x"08", x"0E", x"01", x"F6", x"00", x"FE", x"F5", x"FE", x"0A",
	x"0E", x"03", x"F3", x"F7", x"03", x"11", x"08", x"F5", x"FC", x"00", x"0E", x"FE",
	x"ED", x"F8", x"ED", x"F5", x"FB", x"02", x"16", x"06", x"FE", x"0B", x"05", x"F2",
	x"F1", x"F9", x"01", x"0E", x"05", x"00", x"F3", x"07", x"F9", x"FD", x"06", x"03",
	x"0A", x"07", x"F3", x"F4", x"F4", x"EE", x"F1", x"05", x"12", x"FA", x"FD", x"12",
	x"F6", x"F7", x"0C", x"16", x"00", x"F5", x"FC", x"0D", x"FD", x"FD", x"17", x"0D",
	x"0E", x"07", x"12", x"FD", x"E2", x"F5", x"07", x"0F", x"17", x"0E", x"F4", x"FF",
	x"06", x"09", x"0B", x"FF", x"01", x"1D", x"08", x"FC", x"0D", x"0F", x"0C", x"FA",
	x"0B", x"07", x"F8", x"F8", x"F3", x"0D", x"0E", x"FA", x"E7", x"E7", x"01", x"09",
	x"FD", x"F1", x"E8", x"F2", x"F9", x"FA", x"F3", x"F6", x"F8", x"F1", x"FA", x"F9",
	x"F4", x"F6", x"EE", x"EA", x"F1", x"01", x"0F", x"05", x"FD", x"FD", x"04", x"05",
	x"E6", x"E4", x"FC", x"FE", x"F4", x"EE", x"F0", x"EC", x"F0", x"F7", x"00", x"F7",
	x"E4", x"F1", x"09", x"03", x"F2", x"EA", x"F5", x"F9", x"08", x"18", x"13", x"11",
	x"F0", x"E8", x"F0", x"F2", x"01", x"FE", x"04", x"0D", x"0C", x"FB", x"EF", x"F5",
	x"FC", x"FA", x"00", x"FC", x"F0", x"F1", x"F3", x"08", x"03", x"03", x"05", x"07",
	x"03", x"FA", x"00", x"01", x"06", x"F5", x"F1", x"03", x"00", x"F7", x"01", x"07",
	x"01", x"EF", x"EF", x"05", x"0D", x"0E", x"FC", x"F2", x"FF", x"04", x"12", x"09",
	x"FE", x"0E", x"17", x"12", x"0B", x"10", x"0C", x"0F", x"11", x"00", x"07", x"14",
	x"0D", x"07", x"0D", x"10", x"13", x"08", x"04", x"05", x"01", x"FD", x"03", x"02",
	x"06", x"13", x"11", x"0A", x"03", x"02", x"01", x"06", x"0F", x"15", x"10", x"04",
	x"07", x"0A", x"08", x"F3", x"F6", x"09", x"06", x"04", x"FD", x"EC", x"E9", x"04",
	x"0B", x"F5", x"F4", x"08", x"0F", x"FE", x"FE", x"01", x"FE", x"F7", x"00", x"0B",
	x"09", x"0B", x"08", x"FF", x"01", x"09", x"F6", x"FA", x"03", x"10", x"07", x"F0",
	x"F2", x"EB", x"F0", x"F3", x"0D", x"17", x"0B", x"F1", x"E8", x"05", x"0E", x"0C",
	x"08", x"05", x"F4", x"06", x"01", x"F1", x"EA", x"E6", x"F8", x"F9", x"FA", x"04",
	x"02", x"F7", x"F2", x"F9", x"F8", x"F4", x"ED", x"F8", x"FE", x"F5", x"F5", x"FF",
	x"00", x"FA", x"06", x"08", x"F7", x"E6", x"E3", x"F8", x"07", x"FB", x"F6", x"02",
	x"FF", x"F9", x"EB", x"F3", x"F5", x"F7", x"F4", x"03", x"01", x"EB", x"F8", x"02",
	x"04", x"F5", x"F1", x"F7", x"03", x"02", x"05", x"07", x"03", x"05", x"FD", x"0E",
	x"0A", x"03", x"07", x"10", x"15", x"06", x"07", x"FA", x"00", x"04", x"04", x"0C",
	x"07", x"07", x"05", x"0A", x"06", x"0C", x"0E", x"08", x"06", x"02", x"09", x"14",
	x"23", x"0E", x"00", x"0B", x"1C", x"0A", x"00", x"0C", x"11", x"0C", x"0A", x"0D",
	x"01", x"00", x"04", x"0B", x"0C", x"05", x"F8", x"F1", x"FE", x"02", x"10", x"18",
	x"0C", x"02", x"08", x"02", x"F3", x"00", x"07", x"0A", x"01", x"FA", x"F8", x"F4",
	x"02", x"09", x"FE", x"FF", x"0C", x"0D", x"01", x"F2", x"06", x"0E", x"FB", x"06",
	x"02", x"FD", x"FF", x"FB", x"06", x"07", x"10", x"13", x"00", x"FB", x"04", x"00",
	x"07", x"0C", x"01", x"FF", x"F9", x"FA", x"FD", x"0A", x"0D", x"FA", x"F3", x"EC",
	x"F3", x"00", x"06", x"06", x"0A", x"FE", x"F5", x"FC", x"F8", x"FA", x"09", x"13",
	x"08", x"02", x"05", x"02", x"FD", x"FA", x"FA", x"00", x"04", x"07", x"03", x"FE",
	x"F1", x"F2", x"FF", x"01", x"00", x"FA", x"F9", x"F9", x"F9", x"F6", x"ED", x"F9",
	x"0E", x"02", x"F7", x"F9", x"FA", x"F9", x"F1", x"FA", x"FF", x"00", x"FE", x"08",
	x"07", x"FF", x"FE", x"FD", x"FF", x"FF", x"00", x"F5", x"FA", x"03", x"FD", x"F4",
	x"F2", x"FB", x"0C", x"0C", x"02", x"11", x"10", x"FE", x"ED", x"F0", x"05", x"04",
	x"01", x"01", x"F8", x"F7", x"F8", x"F7", x"0B", x"0E", x"04", x"F9", x"FE", x"FB",
	x"F9", x"F7", x"FF", x"02", x"FE", x"03", x"00", x"FC", x"08", x"FB", x"F9", x"0C",
	x"10", x"0A", x"05", x"02", x"07", x"01", x"0B", x"0E", x"05", x"05", x"00", x"F8",
	x"FA", x"FC", x"FE", x"05", x"09", x"10", x"F9", x"EE", x"F9", x"FF", x"02", x"02",
	x"FE", x"09", x"04", x"FC", x"FC", x"FF", x"07", x"00", x"F7", x"03", x"0A", x"07",
	x"03", x"04", x"0A", x"03", x"FB", x"01", x"07", x"0C", x"FD", x"FB", x"FB", x"F4",
	x"F4", x"04", x"01", x"FC", x"FF", x"F8", x"FB", x"FD", x"FB", x"FA", x"F3", x"F8",
	x"FD", x"01", x"02", x"FA", x"F6", x"01", x"03", x"FD", x"0C", x"0B", x"03", x"FB",
	x"F2", x"FE", x"09", x"09", x"08", x"02", x"FE", x"02", x"0D", x"12", x"12", x"08",
	x"FE", x"F9", x"FD", x"06", x"10", x"11", x"0D", x"0D", x"0F", x"09", x"08", x"09",
	x"06", x"02", x"09", x"0A", x"09", x"03", x"04", x"04", x"F4", x"01", x"09", x"04",
	x"00", x"FE", x"04", x"00", x"05", x"0B", x"07", x"04", x"02", x"11", x"0C", x"03",
	x"06", x"FE", x"03", x"08", x"FF", x"01", x"F5", x"F7", x"06", x"04", x"FF", x"00",
	x"FE", x"F8", x"01", x"06", x"06", x"FF", x"00", x"FD", x"F7", x"FF", x"07", x"07",
	x"03", x"02", x"F5", x"F4", x"FB", x"FC", x"02", x"01", x"F8", x"F2", x"F8", x"FC",
	x"F9", x"FB", x"FB", x"F8", x"FA", x"F4", x"F4", x"F9", x"FE", x"03", x"06", x"F7",
	x"F5", x"FB", x"FF", x"FE", x"F4", x"EC", x"F9", x"F6", x"F3", x"FA", x"FE", x"02",
	x"03", x"FA", x"F8", x"F3", x"F5", x"00", x"FE", x"F8", x"FC", x"05", x"02", x"02",
	x"04", x"FD", x"02", x"00", x"04", x"04", x"04", x"07", x"01", x"F7", x"00", x"0A",
	x"09", x"08", x"09", x"08", x"06", x"FF", x"00", x"05", x"03", x"07", x"0A", x"04",
	x"03", x"0E", x"16", x"14", x"08", x"03", x"FE", x"FE", x"06", x"07", x"0F", x"09",
	x"02", x"05", x"FF", x"06", x"0A", x"09", x"04", x"0B", x"0E", x"0F", x"0B", x"0F",
	x"13", x"08", x"03", x"07", x"09", x"0D", x"0C", x"00", x"05", x"09", x"00", x"FB",
	x"F9", x"FF", x"04", x"03", x"00", x"02", x"02", x"FC", x"FA", x"05", x"04", x"FF",
	x"02", x"06", x"FE", x"EB", x"EE", x"FA", x"05", x"01", x"F4", x"F1", x"F3", x"FC",
	x"F6", x"EF", x"FA", x"FC", x"01", x"FC", x"EC", x"F0", x"F3", x"F9", x"02", x"04",
	x"FC", x"F5", x"F7", x"F8", x"FC", x"01", x"04", x"FD", x"FA", x"FD", x"FA", x"FA",
	x"FD", x"F4", x"F8", x"08", x"03", x"FA", x"F8", x"F7", x"03", x"02", x"F6", x"00",
	x"05", x"FF", x"FD", x"02", x"00", x"F9", x"FC", x"04", x"0A", x"08", x"01", x"F8",
	x"F8", x"FD", x"02", x"05", x"02", x"FE", x"04", x"09", x"0A", x"06", x"FF", x"02",
	x"05", x"06", x"FF", x"F9", x"04", x"0A", x"09", x"0A", x"02", x"04", x"03", x"07",
	x"03", x"02", x"04", x"0D", x"11", x"0C", x"08", x"02", x"FD", x"FF", x"01", x"05",
	x"04", x"03", x"04", x"07", x"04", x"04", x"08", x"00", x"FA", x"FC", x"FF", x"06",
	x"02", x"FF", x"FF", x"FE", x"07", x"0A", x"01", x"FA", x"FB", x"F6", x"F9", x"FF",
	x"FB", x"02", x"FE", x"F9", x"F8", x"F4", x"F8", x"FC", x"F6", x"F4", x"F2", x"F3",
	x"F5", x"FB", x"FA", x"F5", x"F0", x"F4", x"F4", x"F2", x"F8", x"F6", x"F7", x"FD",
	x"FF", x"FA", x"F6", x"FC", x"FC", x"FA", x"00", x"FF", x"F1", x"EA", x"EE", x"FB",
	x"04", x"01", x"FE", x"FA", x"F2", x"F5", x"FC", x"00", x"FD", x"FA", x"03", x"FF",
	x"FA", x"FE", x"FB", x"FE", x"FF", x"01", x"06", x"08", x"08", x"01", x"FE", x"02",
	x"FF", x"03", x"09", x"06", x"06", x"03", x"FB", x"FF", x"08", x"0B", x"09", x"0A",
	x"09", x"0B", x"08", x"09", x"07", x"03", x"02", x"06", x"09", x"0E", x"06", x"05",
	x"07", x"05", x"06", x"09", x"01", x"FE", x"04", x"0D", x"0F", x"0A", x"00", x"F9",
	x"04", x"0C", x"06", x"06", x"FF", x"00", x"02", x"08", x"07", x"FF", x"FF", x"FF",
	x"FA", x"F9", x"FC", x"06", x"06", x"08", x"09", x"FD", x"FB", x"F4", x"F9", x"07",
	x"01", x"FB", x"03", x"01", x"F4", x"F8", x"FC", x"FF", x"02", x"FA", x"FA", x"FE",
	x"F3", x"F1", x"FF", x"FF", x"F8", x"F9", x"FC", x"00", x"00", x"FD", x"FD", x"00",
	x"FE", x"FE", x"01", x"04", x"FF", x"FE", x"01", x"03", x"06", x"04", x"FE", x"F4",
	x"F4", x"FA", x"FE", x"03", x"00", x"01", x"FA", x"FC", x"01", x"00", x"01", x"00",
	x"05", x"01", x"00", x"05", x"00", x"04", x"07", x"06", x"00", x"FF", x"07", x"03",
	x"FE", x"FB", x"03", x"04", x"02", x"FE", x"FB", x"07", x"0A", x"08", x"09", x"08",
	x"08", x"01", x"FF", x"09", x"0D", x"11", x"07", x"FE", x"03", x"06", x"09", x"0B",
	x"02", x"08", x"08", x"06", x"04", x"FD", x"FE", x"02", x"03", x"00", x"FF", x"03",
	x"02", x"00", x"04", x"0B", x"06", x"05", x"04", x"04", x"02", x"02", x"0A", x"04",
	x"FB", x"FF", x"04", x"04", x"03", x"FD", x"FC", x"FD", x"05", x"07", x"02", x"FD",
	x"FB", x"FF", x"08", x"0A", x"03", x"FF", x"FF", x"FF", x"FF", x"FD", x"F8", x"FB",
	x"FD", x"FA", x"FC", x"FC", x"00", x"FD", x"FA", x"00", x"02", x"F9", x"F8", x"FA",
	x"02", x"08", x"01", x"FB", x"FA", x"FA", x"03", x"04", x"01", x"00", x"FD", x"FB",
	x"FA", x"FC", x"FF", x"03", x"00", x"02", x"FE", x"FA", x"FD", x"FB", x"FD", x"03",
	x"08", x"08", x"FC", x"FF", x"05", x"04", x"08", x"05", x"FD", x"FB", x"FE", x"02",
	x"08", x"09", x"02", x"01", x"02", x"06", x"05", x"03", x"0B", x"0D", x"07", x"05",
	x"01", x"06", x"09", x"01", x"FE", x"00", x"06", x"04", x"FF", x"07", x"0A", x"05",
	x"FE", x"FE", x"01", x"FF", x"F9", x"FE", x"01", x"FC", x"FF", x"03", x"01", x"FD",
	x"FD", x"00", x"02", x"01", x"FF", x"FD", x"FD", x"FE", x"00", x"04", x"03", x"0A",
	x"0B", x"03", x"FA", x"F8", x"02", x"0B", x"04", x"02", x"03", x"04", x"02", x"F9",
	x"F6", x"FA", x"01", x"05", x"03", x"FF", x"FB", x"FC", x"FD", x"02", x"03", x"FF",
	x"FE", x"04", x"FF", x"FB", x"FD", x"F9", x"FB", x"F6", x"F6", x"F9", x"FD", x"FD",
	x"00", x"F7", x"EF", x"F5", x"FA", x"03", x"02", x"00", x"FF", x"F9", x"FA", x"01",
	x"FC", x"FD", x"FB", x"FC", x"FF", x"F9", x"F9", x"F7", x"F2", x"F7", x"FA", x"FB",
	x"00", x"FB", x"FE", x"01", x"02", x"FF", x"FE", x"03", x"00", x"00", x"FE", x"00",
	x"FE", x"00", x"06", x"02", x"02", x"03", x"00", x"01", x"05", x"0A", x"0D", x"0D",
	x"0B", x"09", x"04", x"03", x"04", x"04", x"10", x"14", x"0E", x"04", x"FE", x"FE",
	x"03", x"08", x"09", x"07", x"04", x"05", x"07", x"08", x"08", x"03", x"FE", x"05",
	x"0D", x"0B", x"06", x"0B", x"08", x"01", x"07", x"0F", x"0E", x"03", x"00", x"05",
	x"0B", x"0A", x"03", x"00", x"01", x"01", x"03", x"06", x"04", x"03", x"04", x"03",
	x"FB", x"FC", x"00", x"01", x"F8", x"F7", x"00", x"FE", x"FB", x"F4", x"F6", x"FC",
	x"FC", x"FF", x"FB", x"F7", x"F2", x"EF", x"FB", x"04", x"FC", x"F7", x"F8", x"F7",
	x"F9", x"F8", x"F6", x"FC", x"FF", x"FB", x"F5", x"F8", x"F6", x"F5", x"F7", x"FD",
	x"FB", x"F2", x"F3", x"F8", x"F8", x"F4", x"F1", x"F5", x"F8", x"F6", x"F4", x"F3",
	x"F3", x"F4", x"F9", x"F6", x"F4", x"F5", x"FB", x"01", x"FE", x"FA", x"F6", x"FB",
	x"FB", x"F8", x"FA", x"FB", x"00", x"00", x"F9", x"F9", x"FD", x"FD", x"FC", x"FC",
	x"05", x"02", x"FF", x"00", x"01", x"01", x"01", x"03", x"05", x"04", x"03", x"02",
	x"02", x"08", x"0C", x"0A", x"07", x"05", x"0B", x"0D", x"09", x"06", x"07", x"08",
	x"0A", x"0A", x"07", x"06", x"06", x"09", x"0B", x"0E", x"0B", x"09", x"0C", x"0F",
	x"0E", x"0B", x"0D", x"0D", x"0A", x"09", x"08", x"07", x"0A", x"0D", x"0D", x"0F",
	x"09", x"FF", x"00", x"08", x"04", x"04", x"06", x"03", x"04", x"07", x"03", x"03",
	x"05", x"07", x"07", x"00", x"FF", x"03", x"05", x"04", x"FD", x"FC", x"FE", x"00",
	x"03", x"04", x"01", x"FD", x"FC", x"FB", x"F6", x"F9", x"FE", x"00", x"00", x"F8",
	x"F6", x"F6", x"F6", x"F9", x"FF", x"FF", x"FC", x"F7", x"F4", x"F2", x"F4", x"F6",
	x"F4", x"F5", x"F8", x"F6", x"F6", x"FA", x"F9", x"F6", x"F4", x"F6", x"F8", x"F6",
	x"F7", x"FD", x"FD", x"FA", x"F7", x"F6", x"FA", x"FA", x"F4", x"F1", x"F6", x"FA",
	x"FB", x"FA", x"F8", x"F8", x"FF", x"01", x"FC", x"FE", x"02", x"00", x"FF", x"01",
	x"07", x"06", x"01", x"00", x"FF", x"03", x"02", x"00", x"02", x"08", x"07", x"06",
	x"02", x"01", x"FD", x"FF", x"0B", x"0B", x"08", x"04", x"00", x"06", x"05", x"05",
	x"0A", x"0F", x"08", x"04", x"08", x"05", x"06", x"09", x"0B", x"0B", x"09", x"04",
	x"01", x"FE", x"02", x"06", x"06", x"04", x"02", x"03", x"02", x"01", x"FD", x"02",
	x"08", x"07", x"01", x"FE", x"FF", x"04", x"00", x"FE", x"FF", x"05", x"02", x"FF",
	x"FF", x"FC", x"FB", x"FF", x"FF", x"FC", x"F8", x"FB", x"FD", x"FB", x"F7", x"F9",
	x"FB", x"F9", x"FF", x"01", x"FD", x"FB", x"FA", x"F8", x"F8", x"F9", x"FD", x"FC",
	x"FA", x"FD", x"00", x"FE", x"F7", x"F5", x"FA", x"FC", x"FB", x"FC", x"FC", x"FA",
	x"F7", x"F6", x"F7", x"F5", x"F7", x"FB", x"FC", x"FD", x"FB", x"F8", x"FB", x"FF",
	x"FC", x"FE", x"FF", x"01", x"03", x"FF", x"01", x"05", x"01", x"FF", x"FF", x"01",
	x"FF", x"FD", x"FC", x"FF", x"04", x"02", x"FE", x"FB", x"FF", x"05", x"08", x"05",
	x"00", x"01", x"06", x"02", x"01", x"01", x"05", x"06", x"00", x"01", x"03", x"01",
	x"FE", x"02", x"FE", x"FA", x"FA", x"FA", x"FC", x"FD", x"00", x"FF", x"FF", x"00",
	x"FF", x"FE", x"FE", x"02", x"04", x"02", x"02", x"01", x"FF", x"00", x"03", x"07",
	x"06", x"00", x"FE", x"FF", x"FE", x"FE", x"00", x"02", x"02", x"01", x"FE", x"FD",
	x"FE", x"01", x"02", x"00", x"FD", x"FD", x"FB", x"FA", x"FC", x"FD", x"FD", x"FF",
	x"00", x"FA", x"F7", x"F8", x"F8", x"FA", x"FF", x"01", x"01", x"00", x"FC", x"FA",
	x"FA", x"F9", x"FE", x"00", x"FF", x"FC", x"F8", x"F9", x"FA", x"FA", x"F9", x"F7",
	x"FA", x"FD", x"FB", x"F7", x"F9", x"FB", x"FC", x"FD", x"FA", x"F9", x"FF", x"03",
	x"03", x"FF", x"F7", x"F5", x"F8", x"FE", x"01", x"FF", x"FB", x"F8", x"FF", x"02",
	x"FC", x"FA", x"FB", x"00", x"04", x"03", x"01", x"FF", x"00", x"02", x"04", x"03",
	x"03", x"00", x"00", x"01", x"FE", x"FD", x"FC", x"00", x"07", x"04", x"01", x"00",
	x"00", x"00", x"02", x"07", x"02", x"FE", x"FC", x"FD", x"02", x"03", x"02", x"08",
	x"0B", x"04", x"FE", x"FB", x"00", x"03", x"05", x"06", x"01", x"FF", x"FF", x"FF",
	x"FF", x"FD", x"01", x"05", x"03", x"02", x"FB", x"FB", x"FF", x"FE", x"00", x"00",
	x"FD", x"FB", x"FC", x"FF", x"FF", x"00", x"00", x"FC", x"F9", x"FD", x"FE", x"FE",
	x"FA", x"F8", x"FB", x"F9", x"F9", x"F8", x"FB", x"FC", x"F9", x"F9", x"F9", x"FB",
	x"FA", x"FB", x"FB", x"FC", x"FD", x"FC", x"FC", x"FB", x"FC", x"FB", x"FD", x"01",
	x"00", x"FC", x"F7", x"F9", x"FC", x"F9", x"F9", x"F7", x"FB", x"FD", x"FC", x"FD",
	x"FE", x"FF", x"01", x"00", x"FE", x"FE", x"FF", x"FC", x"FE", x"FE", x"FF", x"02",
	x"01", x"FC", x"FA", x"FD", x"FF", x"FE", x"FE", x"FD", x"FE", x"01", x"00", x"01",
	x"03", x"04", x"00", x"FF", x"01", x"00", x"FD", x"FC", x"00", x"05", x"03", x"FF",
	x"FF", x"01", x"05", x"05", x"00", x"00", x"FD", x"00", x"07", x"09", x"07", x"06",
	x"01", x"FF", x"FD", x"FF", x"00", x"01", x"03", x"02", x"02", x"FC", x"FA", x"00",
	x"03", x"01", x"FE", x"FE", x"01", x"02", x"FE", x"01", x"01", x"04", x"06", x"02",
	x"FD", x"FC", x"FD", x"FD", x"00", x"01", x"FD", x"FB", x"FC", x"FF", x"FE", x"FC",
	x"F9", x"FB", x"FF", x"02", x"FF", x"FD", x"FE", x"FE", x"FC", x"FB", x"FE", x"FE",
	x"FC", x"FC", x"FB", x"FA", x"01", x"03", x"FB", x"F3", x"F3", x"FD", x"FF", x"FE",
	x"FB", x"F4", x"F5", x"FA", x"FC", x"FC", x"FA", x"F9", x"FB", x"FC", x"F9", x"F6",
	x"F9", x"FD", x"FD", x"F9", x"FA", x"FF", x"FE", x"F8", x"FA", x"FF", x"FF", x"FA",
	x"F6", x"FA", x"FE", x"FE", x"FB", x"FB", x"00", x"03", x"FE", x"FB", x"FC", x"FE",
	x"FF", x"FF", x"01", x"04", x"00", x"FF", x"FD", x"FD", x"FE", x"FD", x"FE", x"03",
	x"03", x"00", x"01", x"01", x"FF", x"FF", x"01", x"02", x"02", x"00", x"00", x"FF",
	x"02", x"03", x"02", x"03", x"07", x"05", x"01", x"FF", x"00", x"00", x"05", x"05",
	x"01", x"01", x"02", x"03", x"03", x"00", x"FF", x"FE", x"FF", x"01", x"01", x"00",
	x"FD", x"FD", x"00", x"02", x"03", x"FE", x"FB", x"FB", x"FA", x"FC", x"FB", x"FA",
	x"FC", x"FE", x"00", x"FF", x"FE", x"FD", x"FE", x"FD", x"FC", x"FA", x"F9", x"FB",
	x"F9", x"F5", x"F5", x"F9", x"FE", x"FD", x"F8", x"F7", x"F9", x"FE", x"FE", x"F7",
	x"F6", x"FB", x"FF", x"FF", x"FD", x"FE", x"FC", x"FA", x"FA", x"F8", x"F7", x"F8",
	x"F9", x"FB", x"FD", x"FC", x"FC", x"FB", x"F7", x"F8", x"FA", x"FC", x"FE", x"01",
	x"04", x"04", x"02", x"FF", x"FA", x"F8", x"FC", x"00", x"FE", x"FC", x"FB", x"FA",
	x"FA", x"FC", x"FD", x"FD", x"FE", x"FD", x"FE", x"02", x"03", x"01", x"FF", x"FC",
	x"FF", x"02", x"03", x"05", x"01", x"00", x"FF", x"FD", x"FE", x"FE", x"FE", x"04",
	x"08", x"04", x"FF", x"FE", x"00", x"00", x"01", x"02", x"02", x"05", x"07", x"04",
	x"01", x"03", x"04", x"05", x"01", x"FF", x"00", x"02", x"06", x"09", x"06", x"04",
	x"05", x"06", x"03", x"01", x"02", x"03", x"04", x"05", x"07", x"04", x"00", x"03",
	x"08", x"07", x"04", x"03", x"02", x"01", x"01", x"03", x"02", x"01", x"01", x"01",
	x"00", x"FF", x"FF", x"01", x"00", x"FD", x"FE", x"FC", x"FD", x"00", x"01", x"05",
	x"02", x"FE", x"FE", x"F9", x"F9", x"FA", x"FC", x"00", x"02", x"FD", x"FC", x"FB",
	x"F9", x"FB", x"FC", x"FC", x"FD", x"FD", x"FB", x"FB", x"FB", x"FA", x"FA", x"FA",
	x"F8", x"F6", x"F4", x"F6", x"FC", x"00", x"FC", x"F8", x"F8", x"F8", x"F8", x"FA",
	x"FC", x"FF", x"FF", x"FE", x"FB", x"FA", x"FB", x"FE", x"FD", x"FE", x"01", x"FE",
	x"F9", x"F7", x"FA", x"FE", x"01", x"01", x"00", x"FE", x"00", x"01", x"FE", x"FE",
	x"00", x"FE", x"FC", x"FD", x"02", x"03", x"02", x"01", x"05", x"09", x"04", x"FE",
	x"FD", x"00", x"02", x"02", x"03", x"03", x"01", x"01", x"03", x"07", x"07", x"01",
	x"02", x"06", x"05", x"01", x"FD", x"00", x"05", x"05", x"05", x"06", x"05", x"02",
	x"02", x"05", x"05", x"06", x"05", x"01", x"00", x"01", x"01", x"01", x"03", x"07",
	x"05", x"00", x"FE", x"01", x"02", x"00", x"FE", x"FF", x"03", x"05", x"03", x"01",
	x"FD", x"00", x"01", x"FF", x"FF", x"FF", x"FE", x"FE", x"00", x"FD", x"FA", x"00",
	x"00", x"FC", x"FE", x"FE", x"FE", x"FF", x"FE", x"FB", x"FA", x"FC", x"FB", x"F8",
	x"FE", x"00", x"FE", x"FE", x"FF", x"FE", x"FF", x"02", x"00", x"01", x"04", x"02",
	x"FE", x"FD", x"FF", x"00", x"FE", x"FF", x"FE", x"FB", x"FD", x"FF", x"00", x"FD",
	x"FF", x"00", x"FE", x"FC", x"FD", x"00", x"04", x"08", x"07", x"03", x"FE", x"FC",
	x"FF", x"03", x"05", x"00", x"FE", x"01", x"00", x"FC", x"00", x"06", x"04", x"00",
	x"FF", x"05", x"06", x"02", x"FE", x"FC", x"01", x"01", x"FE", x"FD", x"FF", x"00",
	x"01", x"05", x"04", x"FF", x"FC", x"FC", x"FD", x"01", x"01", x"FE", x"FD", x"00",
	x"00", x"FF", x"00", x"01", x"FF", x"FD", x"FC", x"FB", x"FE", x"FE", x"FD", x"00",
	x"00", x"00", x"03", x"02", x"FF", x"FC", x"FE", x"FF", x"FD", x"FC", x"FC", x"FD",
	x"FB", x"F9", x"FB", x"FE", x"FD", x"FB", x"FB", x"FC", x"FA", x"F9", x"FE", x"00",
	x"FC", x"F9", x"F6", x"F8", x"F9", x"F9", x"FB", x"FD", x"FD", x"FA", x"F9", x"FA",
	x"FB", x"FC", x"FD", x"FE", x"FD", x"F9", x"F8", x"FC", x"FF", x"FE", x"FB", x"F9",
	x"FC", x"FC", x"FD", x"FE", x"FE", x"FE", x"FC", x"FD", x"FC", x"FE", x"00", x"02",
	x"02", x"FE", x"00", x"04", x"02", x"FF", x"01", x"02", x"01", x"01", x"FE", x"FF",
	x"FF", x"FE", x"FD", x"FF", x"03", x"03", x"02", x"00", x"02", x"05", x"04", x"04",
	x"04", x"04", x"02", x"01", x"00", x"01", x"03", x"03", x"01", x"02", x"04", x"02",
	x"02", x"05", x"05", x"03", x"01", x"00", x"FF", x"FF", x"01", x"02", x"02", x"04",
	x"03", x"FF", x"FF", x"01", x"01", x"FF", x"00", x"FE", x"FA", x"FA", x"FD", x"FF",
	x"FF", x"00", x"00", x"FF", x"FE", x"FD", x"FB", x"FC", x"FD", x"FF", x"FE", x"FF",
	x"FE", x"FD", x"FC", x"FC", x"FD", x"00", x"01", x"FE", x"FB", x"FB", x"FD", x"00",
	x"FF", x"FF", x"FD", x"FC", x"FF", x"00", x"FE", x"FE", x"FF", x"FF", x"00", x"FF",
	x"00", x"FE", x"FE", x"00", x"FF", x"FD", x"00", x"02", x"01", x"00", x"00", x"01",
	x"FF", x"FE", x"02", x"05", x"03", x"FE", x"FF", x"01", x"01", x"00", x"00", x"02",
	x"04", x"05", x"00", x"FD", x"FE", x"00", x"02", x"02", x"02", x"02", x"03", x"FF",
	x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"FE", x"FD", x"FE", x"FF", x"FE", x"FC",
	x"FC", x"FF", x"00", x"FF", x"FD", x"FD", x"00", x"00", x"00", x"FE", x"FA", x"FC",
	x"00", x"00", x"FC", x"FB", x"FB", x"F9", x"F7", x"F7", x"F9", x"FD", x"FE", x"01",
	x"01", x"FB", x"F8", x"FB", x"00", x"FF", x"FD", x"FE", x"FB", x"FB", x"FB", x"FB",
	x"FC", x"FB", x"FC", x"FE", x"FF", x"FF", x"FB", x"FA", x"FD", x"FD", x"FD", x"FF",
	x"FF", x"FD", x"FD", x"00", x"03", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"02",
	x"01", x"FD", x"FE", x"FF", x"FF", x"00", x"FE", x"00", x"02", x"02", x"00", x"FF",
	x"00", x"01", x"01", x"01", x"02", x"02", x"00", x"FF", x"FF", x"02", x"01", x"FF",
	x"02", x"03", x"FF", x"FF", x"02", x"04", x"05", x"05", x"06", x"05", x"03", x"03",
	x"05", x"04", x"02", x"01", x"02", x"04", x"02", x"FF", x"FF", x"01", x"03", x"02",
	x"01", x"00", x"FE", x"FE", x"02", x"03", x"01", x"FE", x"FF", x"01", x"00", x"00",
	x"00", x"00", x"01", x"02", x"02", x"00", x"FF", x"FF", x"00", x"FF", x"FC", x"FE",
	x"FF", x"FD", x"FE", x"00", x"FF", x"FF", x"FE", x"FE", x"FB", x"FA", x"FE", x"FE",
	x"FC", x"FD", x"00", x"FF", x"00", x"FE", x"FD", x"FE", x"FC", x"FD", x"FF", x"00",
	x"FF", x"FE", x"FD", x"FC", x"FC", x"FE", x"FF", x"FF", x"FD", x"FD", x"FF", x"FD",
	x"FA", x"FB", x"FF", x"01", x"FD", x"FE", x"02", x"FF", x"FA", x"F8", x"FB", x"FF",
	x"00", x"01", x"00", x"FF", x"FD", x"F9", x"FB", x"FB", x"FD", x"00", x"FF", x"FD",
	x"FC", x"FD", x"FE", x"FE", x"FE", x"FB", x"FB", x"FE", x"01", x"00", x"FD", x"FE",
	x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FE",
	x"FC", x"FD", x"FF", x"FE", x"FD", x"00", x"02", x"01", x"FE", x"FF", x"00", x"FE",
	x"FE", x"FF", x"02", x"02", x"02", x"01", x"02", x"01", x"01", x"03", x"04", x"04",
	x"01", x"01", x"02", x"01", x"02", x"01", x"02", x"02", x"03", x"02", x"01", x"01",
	x"01", x"02", x"02", x"02", x"03", x"03", x"02", x"03", x"02", x"02", x"03", x"03",
	x"04", x"02", x"01", x"02", x"03", x"03", x"03", x"02", x"00", x"FF", x"FE", x"FE",
	x"00", x"01", x"01", x"FF", x"00", x"00", x"02", x"03", x"02", x"00", x"FE", x"FF",
	x"FF", x"FF", x"FC", x"FD", x"FF", x"FF", x"FE", x"FF", x"FD", x"FC", x"FD", x"FE",
	x"FD", x"FC", x"FD", x"FD", x"FC", x"FB", x"FC", x"FC", x"FC", x"FC", x"FA", x"FB",
	x"FB", x"FA", x"FB", x"FA", x"FA", x"FC", x"FF", x"FE", x"FB", x"FA", x"FC", x"FB",
	x"FC", x"FC", x"FA", x"FA", x"FB", x"FC", x"FF", x"FE", x"FD", x"FC", x"FE", x"FF",
	x"FD", x"FC", x"FC", x"FD", x"00", x"00", x"FE", x"FE", x"01", x"02", x"00", x"FF",
	x"FF", x"FE", x"02", x"02", x"01", x"01", x"02", x"03", x"00", x"00", x"02", x"03",
	x"01", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"03", x"03", x"04",
	x"05", x"04", x"05", x"03", x"01", x"01", x"02", x"04", x"05", x"03", x"02", x"02",
	x"04", x"06", x"04", x"02", x"01", x"02", x"05", x"05", x"01", x"FD", x"FE", x"00",
	x"01", x"00", x"00", x"03", x"01", x"FE", x"FE", x"FE", x"FE", x"FC", x"FE", x"00",
	x"FF", x"FE", x"FB", x"FC", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FD",
	x"FD", x"FC", x"FD", x"FE", x"FF", x"FE", x"FB", x"FB", x"FF", x"FF", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FE", x"FD", x"FD", x"FE", x"FD", x"FB", x"FD", x"FF", x"FD",
	x"FD", x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"01", x"02", x"00", x"FD", x"FD",
	x"FF", x"01", x"01", x"FF", x"FD", x"FF", x"00", x"01", x"00", x"01", x"01", x"01",
	x"00", x"00", x"00", x"FF", x"00", x"03", x"05", x"04", x"04", x"04", x"01", x"00",
	x"03", x"04", x"01", x"01", x"02", x"02", x"00", x"00", x"02", x"04", x"02", x"00",
	x"01", x"02", x"02", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"02",
	x"01", x"02", x"00", x"FF", x"00", x"03", x"03", x"01", x"00", x"00", x"02", x"03",
	x"00", x"FF", x"00", x"00", x"01", x"00", x"01", x"00", x"FF", x"01", x"02", x"03",
	x"02", x"FF", x"FD", x"FD", x"FE", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FD", x"FC", x"FF", x"FF", x"FC", x"FB", x"FD", x"01", x"02", x"00", x"FF",
	x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"01", x"03", x"00", x"FD", x"FD", x"FE", x"FE", x"FF", x"01", x"01", x"FD", x"FB",
	x"FD", x"FE", x"FE", x"FF", x"01", x"01", x"FF", x"FD", x"FE", x"FE", x"FE", x"FF",
	x"00", x"03", x"02", x"FF", x"FE", x"01", x"03", x"02", x"00", x"FF", x"00", x"FF",
	x"FF", x"00", x"FF", x"00", x"01", x"00", x"00", x"01", x"01", x"00", x"00", x"01",
	x"00", x"FF", x"FF", x"01", x"02", x"03", x"03", x"00", x"FE", x"00", x"03", x"04",
	x"03", x"03", x"02", x"00", x"FF", x"FF", x"FF", x"01", x"02", x"03", x"04", x"03",
	x"01", x"00", x"02", x"03", x"FF", x"FF", x"00", x"01", x"FF", x"00", x"03", x"04",
	x"02", x"00", x"01", x"02", x"00", x"00", x"02", x"03", x"04", x"04", x"03", x"01",
	x"01", x"02", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"01", x"02", x"01",
	x"01", x"01", x"FE", x"FB", x"FD", x"00", x"01", x"FF", x"FD", x"FE", x"FF", x"FE",
	x"FD", x"FE", x"FF", x"FE", x"FC", x"FC", x"FD", x"FE", x"FD", x"FD", x"FE", x"FF",
	x"00", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"FE", x"FF", x"00", x"01", x"01",
	x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"01", x"00", x"FE",
	x"FE", x"FE", x"FF", x"01", x"01", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"02",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"FF", x"FE",
	x"FE", x"00", x"01", x"01", x"FF", x"FD", x"FF", x"00", x"00", x"02", x"03", x"01",
	x"00", x"00", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"01", x"01",
	x"00", x"01", x"02", x"FF", x"FE", x"FE", x"FE", x"00", x"00", x"FF", x"FE", x"FF",
	x"00", x"FF", x"FD", x"FD", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"FF", x"FE", x"FE", x"00", x"00", x"01", x"01", x"00", x"FE", x"FD", x"FD", x"FE",
	x"FE", x"00", x"00", x"00", x"FF", x"FD", x"FE", x"FF", x"FE", x"FE", x"FF", x"00",
	x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE",
	x"00", x"FF", x"FD", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"01", x"02", x"02", x"02", x"03", x"01", x"00", x"00", x"01", x"02", x"03", x"03",
	x"03", x"02", x"02", x"02", x"02", x"02", x"03", x"02", x"02", x"01", x"01", x"00",
	x"FF", x"01", x"01", x"01", x"00", x"FF", x"00", x"01", x"00", x"FF", x"00", x"01",
	x"02", x"02", x"01", x"01", x"00", x"00", x"FF", x"01", x"FF", x"FD", x"FD", x"FE",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"01",
	x"FF", x"FD", x"FF", x"00", x"FF", x"FE", x"00", x"FE", x"FC", x"FC", x"FD", x"00",
	x"00", x"FD", x"FC", x"FC", x"FF", x"FF", x"FD", x"FE", x"FF", x"FE", x"FE", x"FE",
	x"00", x"00", x"FF", x"FF", x"00", x"FE", x"FD", x"FD", x"FE", x"FE", x"00", x"00",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FC", x"FC",
	x"FF", x"00", x"FF", x"FD", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"00", x"FD", x"FD", x"FE", x"FF", x"FF",
	x"02", x"03", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"02", x"01",
	x"FF", x"FE", x"FF", x"FF", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"00", x"01", x"01", x"01", x"FF", x"FF", x"01", x"01", x"00", x"FC",
	x"FD", x"FF", x"02", x"02", x"01", x"FF", x"00", x"02", x"02", x"02", x"01", x"FF",
	x"FE", x"FE", x"00", x"01", x"00", x"01", x"00", x"FF", x"FE", x"FE", x"00", x"00",
	x"00", x"00", x"01", x"01", x"FF", x"00", x"02", x"04", x"02", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"01", x"02", x"02", x"00", x"00", x"00", x"02", x"02", x"00", x"FF", x"FE", x"FF",
	x"00", x"00", x"00", x"00", x"01", x"01", x"FF", x"FD", x"FD", x"FF", x"00", x"00",
	x"FF", x"FE", x"FE", x"FD", x"FF", x"00", x"00", x"01", x"00", x"FE", x"FE", x"01",
	x"02", x"01", x"00", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FE", x"FE", x"FE", x"00", x"01", x"01", x"00", x"FF", x"FD", x"FE", x"FE", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"FF", x"FE", x"FD", x"FD",
	x"FC", x"FD", x"FF", x"FF", x"FE", x"FC", x"FB", x"FC", x"FD", x"FF", x"FE", x"FD",
	x"FC", x"FD", x"FD", x"FC", x"FD", x"00", x"01", x"00", x"FE", x"FD", x"FD", x"FD",
	x"FD", x"FE", x"00", x"FF", x"FC", x"FC", x"FD", x"FF", x"00", x"00", x"FF", x"FE",
	x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"FD", x"FB", x"FC", x"FE",
	x"00", x"01", x"FF", x"FE", x"FF", x"00", x"00", x"01", x"02", x"02", x"00", x"FF",
	x"FF", x"FF", x"01", x"02", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"01", x"01",
	x"00", x"00", x"FF", x"00", x"02", x"03", x"02", x"03", x"04", x"03", x"02", x"01",
	x"03", x"04", x"04", x"03", x"02", x"00", x"FF", x"00", x"02", x"03", x"02", x"02",
	x"01", x"02", x"02", x"01", x"00", x"00", x"02", x"03", x"03", x"01", x"00", x"FF",
	x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"FF", x"FE", x"FD", x"FF",
	x"00", x"FF", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"FE", x"FD", x"FC", x"FC",
	x"FD", x"FD", x"FE", x"FE", x"FF", x"FE", x"FD", x"FC", x"FB", x"FD", x"FE", x"FE",
	x"FC", x"FC", x"FD", x"FE", x"00", x"00", x"FF", x"FD", x"FD", x"FE", x"FF", x"00",
	x"FF", x"FD", x"FD", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE",
	x"FD", x"FC", x"FC", x"FE", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"00", x"00",
	x"00", x"00", x"02", x"02", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"03",
	x"04", x"02", x"FF", x"FF", x"01", x"04", x"04", x"03", x"01", x"00", x"00", x"00",
	x"00", x"00", x"01", x"01", x"00", x"00", x"01", x"02", x"03", x"03", x"03", x"04",
	x"02", x"00", x"FF", x"FF", x"01", x"03", x"02", x"00", x"FF", x"00", x"01", x"00",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"00", x"FF", x"00", x"02", x"02", x"FF",
	x"FE", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"02", x"02", x"01", x"FF",
	x"FF", x"00", x"01", x"01", x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"02", x"02",
	x"01", x"01", x"01", x"00", x"FF", x"FF", x"00", x"01", x"FF", x"FF", x"00", x"00",
	x"01", x"01", x"01", x"00", x"00", x"00", x"01", x"02", x"03", x"02", x"01", x"02",
	x"03", x"02", x"01", x"01", x"02", x"03", x"03", x"01", x"00", x"00", x"00", x"03",
	x"04", x"03", x"01", x"00", x"01", x"02", x"02", x"02", x"01", x"01", x"02", x"02",
	x"01", x"01", x"01", x"02", x"02", x"02", x"02", x"01", x"01", x"01", x"01", x"01",
	x"01", x"00", x"01", x"01", x"01", x"00", x"FE", x"FE", x"FF", x"00", x"00", x"FF",
	x"00", x"02", x"02", x"00", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"FF",
	x"00", x"00", x"00", x"01", x"01", x"01", x"FF", x"FE", x"FF", x"00", x"00", x"FF",
	x"00", x"01", x"00", x"FF", x"FE", x"FF", x"00", x"02", x"01", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FE", x"FF", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FF",
	x"00", x"00", x"FF", x"FD", x"FD", x"FE", x"00", x"00", x"FE", x"FE", x"00", x"02",
	x"01", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"01",
	x"00", x"FE", x"FF", x"01", x"02", x"02", x"01", x"01", x"02", x"02", x"02", x"01",
	x"00", x"00", x"02", x"03", x"03", x"01", x"01", x"03", x"02", x"02", x"03", x"03",
	x"02", x"00", x"00", x"01", x"01", x"02", x"03", x"02", x"02", x"01", x"02", x"02",
	x"01", x"01", x"00", x"01", x"02", x"01", x"01", x"00", x"00", x"00", x"00", x"01",
	x"01", x"01", x"01", x"00", x"FE", x"FE", x"00", x"01", x"00", x"FF", x"FE", x"FD",
	x"FE", x"FE", x"FE", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FD", x"FD", x"FF",
	x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FD", x"FD", x"FE", x"FD", x"FE",
	x"00", x"FF", x"FE", x"FD", x"FE", x"FE", x"FD", x"FD", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"02", x"01", x"01", x"00", x"FF", x"FF", x"01", x"01", x"00", x"00", x"01",
	x"01", x"00", x"00", x"00", x"00", x"01", x"01", x"02", x"01", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"FE", x"FD", x"FF", x"FF",
	x"FF", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FF", x"FE", x"FE", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"00",
	x"01", x"00", x"00", x"FF", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"00",
	x"01", x"00", x"FF", x"01", x"02", x"01", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"01", x"00", x"01", x"02", x"02", x"01", x"01", x"02", x"02", x"02",
	x"03", x"03", x"02", x"02", x"02", x"03", x"03", x"02", x"01", x"01", x"01", x"02",
	x"02", x"02", x"02", x"01", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"01", x"00",
	x"FF", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"00", x"00",
	x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01",
	x"FF", x"FE", x"00", x"01", x"02", x"01", x"01", x"01", x"00", x"00", x"01", x"01",
	x"01", x"01", x"01", x"01", x"00", x"01", x"02", x"01", x"01", x"00", x"00", x"00",
	x"00", x"01", x"01", x"01", x"01", x"02", x"02", x"01", x"00", x"00", x"01", x"02",
	x"02", x"02", x"01", x"01", x"01", x"01", x"02", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"00", x"01", x"02", x"02", x"01", x"01", x"01", x"01", x"01", x"02",
	x"01", x"FF", x"FF", x"00", x"02", x"03", x"02", x"01", x"00", x"00", x"00", x"01",
	x"01", x"01", x"01", x"01", x"02", x"01", x"00", x"00", x"01", x"01", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"02", x"02", x"01", x"00", x"00", x"01", x"02", x"02", x"01", x"00", x"FF", x"00",
	x"00", x"01", x"01", x"01", x"00", x"FE", x"FE", x"FF", x"FE", x"FE", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"01",
	x"FF", x"FE", x"FD", x"FE", x"00", x"01", x"01", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"FF", x"00", x"01", x"01", x"01", x"00", x"01", x"01", x"01", x"01", x"01",
	x"01", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FE", x"FE", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE",
	x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FD", x"FD", x"FC", x"FB", x"FB", x"FC",
	x"FC", x"FC", x"FD", x"FF", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"FE",
	x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"FD", x"FE", x"FF", x"00", x"FF",
	x"FE", x"FE", x"FE", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"00",
	x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01",
	x"01", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00",
	x"01", x"01", x"00", x"FF", x"FF", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"00",
	x"01", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FE", x"FF",
	x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FC", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FD",
	x"FD", x"FE", x"FE", x"FD", x"FC", x"FC", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE", x"FF", x"00", x"FF", x"FF", x"FE",
	x"FD", x"FC", x"FD", x"FE", x"FE", x"FE", x"FE", x"FF", x"FE", x"FE", x"FF", x"00",
	x"00", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"FF",
	x"FE", x"FE", x"FF", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"01", x"01", x"00", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FE", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FE", x"FD", x"FC", x"FC", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FC", x"FC", x"FD", x"FD", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FD", x"FE", x"FE", x"FE", x"FD", x"FC", x"FD", x"FE", x"FE", x"FD", x"FD", x"FD",
	x"FE", x"FE", x"FF", x"FF", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"00", x"00", x"01", x"01", x"02", x"01", x"00", x"00",
	x"01", x"02", x"01", x"00", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"01", x"01",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"00", x"FF", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"FE", x"FF", x"00", x"FF", x"FE", x"FE", x"FD", x"FD",
	x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"01", x"01", x"00",
	x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"01", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"00", x"01", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"FF", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"01", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"01", x"02", x"01", x"01", x"00", x"01", x"01", x"00", x"00", x"00",
	x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"01", x"01", x"01", x"01", x"01",
	x"01", x"00", x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"FE", x"FD",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FE",
	x"FF", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FD",
	x"FD", x"FF", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"01", x"01",
	x"02", x"01", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"01", x"01", x"01", x"00", x"01", x"01", x"01", x"02",
	x"01", x"01", x"00", x"FF", x"FF", x"00", x"01", x"01", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"01",
	x"01", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"01",
	x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00",
	x"FF", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"01", x"01", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"00",
	x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"01",
	x"01", x"00", x"FF", x"FF", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"01", x"02", x"02", x"02", x"01", x"01", x"00", x"00", x"01", x"02", x"02",
	x"01", x"01", x"01", x"01", x"01", x"01", x"02", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"01", x"01", x"02",
	x"02", x"02", x"01", x"01", x"01", x"00", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01"
);

	
signal cnt_out: integer := 0;	
signal play_sound: std_logic := '0';
constant cnt_max: integer := 8857;
--signal out_signal: signed(7 downto 0) := x"00";

begin
	
process (CLK)
begin
    if rising_edge(CLK) then
        if RST = '1' then
            play_sound <= '0';
        elsif PLAY = '1' then
            play_sound <= '1';
        elsif PLAY = '0' and cnt_out = cnt_max then
            play_sound <= '0';
        end if;
    end if;
end process;

	
-- 12bit counter
process (CLK)
begin     
    if rising_edge(CLK) then
        if RST = '1' then
            cnt_out <= 0;
        elsif CE = '1' and play_sound = '1' then
            cnt_out <= cnt_out + 1;       
        end if;
        if cnt_out = cnt_max then
            cnt_out <= 0;            
        end if;        
    end if;
end process;

--SAMPLE_OUT <= kick_sound(conv_integer(cnt_out));
process (CLK) 
begin
    if rising_edge(CLK) then
        if RST = '1' then
            SAMPLE_OUT <= x"00";
        elsif CE = '1' then
            SAMPLE_OUT <= hhat_sound(cnt_out);
        end if;
    end if;    
end process;


end Behavioral;