----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 25.12.2018 17:39:59
-- Design Name: 
-- Module Name: Crash - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Crash is
    Port ( CLK : in STD_LOGIC;
           CE : in STD_LOGIC;
           RST : in STD_LOGIC;
           PLAY : in STD_LOGIC;
           SAMPLE_OUT : out signed(7 downto 0)
           );
end Crash;

architecture Behavioral of Crash is

type memory is array (0 to 18687) of signed(7 downto 0);
constant crash_sound: memory := (
	x"01", x"02", x"FE", x"FD", x"FF", x"09", x"FE", x"FC", x"F6", x"FF", x"06", x"09",
	x"FF", x"FF", x"05", x"07", x"F9", x"F4", x"F3", x"FE", x"FF", x"02", x"06", x"0E",
	x"0D", x"01", x"F9", x"F7", x"F6", x"FB", x"F9", x"FB", x"00", x"12", x"08", x"FF",
	x"FA", x"02", x"03", x"00", x"ED", x"EE", x"FD", x"11", x"11", x"10", x"03", x"F8",
	x"F6", x"F1", x"F1", x"FB", x"09", x"FD", x"FE", x"14", x"14", x"07", x"FA", x"EC",
	x"F6", x"00", x"FE", x"F9", x"FA", x"05", x"FD", x"08", x"04", x"05", x"04", x"04",
	x"01", x"FA", x"FA", x"F4", x"F8", x"05", x"FD", x"01", x"05", x"04", x"0A", x"00",
	x"02", x"F6", x"FE", x"FD", x"FA", x"FC", x"04", x"F7", x"0A", x"02", x"F6", x"FA",
	x"04", x"07", x"0E", x"0C", x"FF", x"F7", x"F7", x"F9", x"F7", x"F0", x"F0", x"02",
	x"08", x"0F", x"10", x"0F", x"0C", x"00", x"F3", x"F9", x"F3", x"F8", x"F4", x"F7",
	x"01", x"FC", x"01", x"08", x"1D", x"11", x"EB", x"F5", x"F1", x"04", x"11", x"0C",
	x"FD", x"F2", x"FE", x"00", x"F3", x"F9", x"FA", x"08", x"02", x"04", x"01", x"FC",
	x"07", x"0D", x"04", x"F3", x"F7", x"FC", x"FB", x"FE", x"0C", x"FE", x"01", x"F8",
	x"FF", x"01", x"0A", x"F9", x"EF", x"08", x"0E", x"FD", x"FB", x"F7", x"0C", x"FB",
	x"0B", x"F8", x"FA", x"FF", x"0E", x"F8", x"00", x"F3", x"01", x"FF", x"02", x"FC",
	x"0F", x"02", x"02", x"F8", x"FE", x"FD", x"03", x"FF", x"FA", x"04", x"11", x"FC",
	x"FB", x"F2", x"FB", x"FF", x"14", x"F7", x"F7", x"FA", x"08", x"F4", x"06", x"05",
	x"0F", x"03", x"06", x"F2", x"F5", x"ED", x"06", x"FE", x"01", x"17", x"0F", x"02",
	x"07", x"EB", x"EC", x"F9", x"ED", x"00", x"FE", x"0E", x"0D", x"16", x"0A", x"FB",
	x"FD", x"FE", x"E9", x"F0", x"0D", x"F6", x"ED", x"0D", x"02", x"0B", x"F6", x"06",
	x"13", x"13", x"08", x"F2", x"EC", x"F7", x"F9", x"FE", x"E0", x"FB", x"11", x"09",
	x"0F", x"14", x"FA", x"0B", x"09", x"F5", x"D6", x"F7", x"05", x"F8", x"FB", x"1E",
	x"08", x"0D", x"FB", x"F1", x"F5", x"08", x"0E", x"FA", x"F6", x"FF", x"06", x"0C",
	x"F7", x"EB", x"E2", x"11", x"FC", x"07", x"03", x"28", x"0C", x"01", x"EB", x"02",
	x"E6", x"05", x"E5", x"FB", x"FF", x"17", x"1E", x"0A", x"E8", x"08", x"F7", x"F9",
	x"EE", x"E6", x"04", x"21", x"0A", x"08", x"FA", x"10", x"F9", x"F5", x"F7", x"EA",
	x"F0", x"1E", x"01", x"F9", x"0A", x"12", x"FE", x"FA", x"0A", x"E3", x"F0", x"02",
	x"FF", x"08", x"04", x"0D", x"05", x"00", x"02", x"F3", x"11", x"F8", x"E8", x"E8",
	x"03", x"0A", x"18", x"02", x"06", x"EE", x"0B", x"EA", x"F7", x"03", x"06", x"14",
	x"14", x"03", x"EF", x"F9", x"00", x"F3", x"E3", x"F7", x"06", x"0F", x"23", x"06",
	x"F5", x"03", x"0D", x"E4", x"DA", x"FB", x"11", x"03", x"0D", x"09", x"F7", x"02",
	x"05", x"FA", x"F6", x"FD", x"15", x"0A", x"ED", x"04", x"F0", x"02", x"03", x"FC",
	x"E4", x"14", x"21", x"05", x"DA", x"03", x"26", x"FC", x"D9", x"DE", x"F4", x"07",
	x"18", x"0E", x"06", x"1F", x"11", x"EF", x"E1", x"F7", x"08", x"FA", x"08", x"FB",
	x"F2", x"0A", x"19", x"EE", x"E4", x"02", x"16", x"04", x"F1", x"FF", x"1A", x"F9",
	x"EC", x"E0", x"FB", x"18", x"2E", x"F3", x"08", x"FC", x"14", x"E7", x"EB", x"EE",
	x"FF", x"06", x"02", x"F3", x"01", x"0F", x"2E", x"F1", x"DD", x"12", x"21", x"F5",
	x"EF", x"DE", x"FD", x"0D", x"01", x"E8", x"F7", x"29", x"1C", x"ED", x"E2", x"0B",
	x"01", x"01", x"F0", x"0E", x"07", x"22", x"07", x"ED", x"DE", x"05", x"01", x"F1",
	x"E1", x"09", x"0C", x"1F", x"0B", x"F5", x"F7", x"04", x"11", x"CE", x"F0", x"19",
	x"14", x"0A", x"06", x"FE", x"F9", x"0E", x"F6", x"F1", x"D7", x"1E", x"F1", x"0C",
	x"06", x"18", x"12", x"F1", x"EC", x"D9", x"FF", x"02", x"09", x"F2", x"09", x"35",
	x"0F", x"EA", x"F2", x"F4", x"F2", x"0E", x"04", x"F6", x"02", x"16", x"F9", x"F2",
	x"07", x"07", x"08", x"EA", x"DF", x"FA", x"03", x"13", x"FD", x"03", x"1D", x"1B",
	x"01", x"D7", x"E6", x"0C", x"14", x"DF", x"FF", x"FE", x"24", x"EE", x"03", x"ED",
	x"04", x"10", x"F0", x"F5", x"03", x"21", x"17", x"F1", x"00", x"F2", x"E9", x"EC",
	x"08", x"E8", x"1D", x"24", x"19", x"E4", x"E6", x"04", x"08", x"E5", x"E9", x"FD",
	x"10", x"1F", x"14", x"F3", x"FA", x"F4", x"0B", x"FC", x"06", x"FD", x"03", x"06",
	x"03", x"E6", x"E7", x"02", x"1C", x"0D", x"DB", x"07", x"11", x"F7", x"FD", x"F8",
	x"0B", x"14", x"19", x"E6", x"DB", x"FC", x"09", x"0A", x"0A", x"F9", x"F3", x"16",
	x"1B", x"E2", x"DC", x"0C", x"28", x"F2", x"E0", x"E2", x"24", x"13", x"03", x"FE",
	x"F8", x"06", x"00", x"06", x"DE", x"F9", x"11", x"1A", x"F1", x"F8", x"EB", x"1D",
	x"12", x"FB", x"D6", x"06", x"2A", x"01", x"D1", x"F5", x"02", x"0E", x"FE", x"F6",
	x"FD", x"1B", x"29", x"00", x"E7", x"01", x"FE", x"F2", x"EF", x"F8", x"EB", x"1B",
	x"13", x"FE", x"CE", x"10", x"03", x"17", x"FA", x"FD", x"0C", x"25", x"0C", x"F7",
	x"F3", x"F5", x"ED", x"FD", x"D8", x"E4", x"07", x"19", x"13", x"16", x"02", x"11",
	x"06", x"01", x"CC", x"ED", x"16", x"07", x"03", x"0E", x"F1", x"02", x"03", x"F9",
	x"EA", x"03", x"11", x"F3", x"0E", x"03", x"F6", x"2B", x"08", x"E0", x"D5", x"02",
	x"F8", x"0C", x"F6", x"F7", x"0F", x"21", x"07", x"ED", x"0E", x"FD", x"F3", x"FE",
	x"EA", x"E6", x"1B", x"0D", x"1B", x"08", x"0B", x"EE", x"F5", x"F5", x"DE", x"EE",
	x"14", x"12", x"0D", x"06", x"FE", x"FB", x"FE", x"E4", x"E1", x"04", x"18", x"24",
	x"2E", x"01", x"EF", x"D6", x"F9", x"F1", x"EE", x"F2", x"12", x"1E", x"18", x"F5",
	x"01", x"03", x"05", x"DA", x"E2", x"F5", x"32", x"14", x"F4", x"F2", x"19", x"16",
	x"E6", x"DC", x"E5", x"04", x"1A", x"08", x"FC", x"EA", x"19", x"2D", x"00", x"D7",
	x"0A", x"01", x"0C", x"EC", x"F8", x"EE", x"1B", x"11", x"D9", x"D5", x"15", x"0D",
	x"07", x"FE", x"FC", x"1D", x"25", x"EA", x"ED", x"E8", x"0D", x"15", x"EF", x"E7",
	x"FF", x"1C", x"03", x"EE", x"F9", x"FE", x"15", x"23", x"E9", x"D7", x"07", x"05",
	x"FB", x"F7", x"03", x"17", x"1B", x"F0", x"E5", x"EE", x"14", x"0A", x"F1", x"EA",
	x"02", x"33", x"11", x"F0", x"0A", x"05", x"F1", x"F0", x"DC", x"DC", x"FA", x"29",
	x"0B", x"FE", x"0B", x"1D", x"F4", x"05", x"EF", x"F2", x"09", x"FD", x"EC", x"FC",
	x"15", x"0D", x"14", x"F2", x"F7", x"F5", x"F2", x"F2", x"01", x"F8", x"25", x"20",
	x"F7", x"E3", x"0A", x"27", x"D7", x"EA", x"EA", x"06", x"07", x"13", x"FD", x"F8",
	x"01", x"0B", x"E1", x"09", x"0A", x"0F", x"07", x"F6", x"13", x"FC", x"1E", x"FB",
	x"DD", x"D7", x"FA", x"0E", x"F7", x"F3", x"32", x"FF", x"EB", x"F9", x"0F", x"09",
	x"EE", x"05", x"E5", x"1D", x"2C", x"F4", x"D7", x"06", x"04", x"E8", x"02", x"F8",
	x"FC", x"0A", x"31", x"FB", x"03", x"E7", x"06", x"03", x"EF", x"E1", x"05", x"08",
	x"0A", x"FA", x"F6", x"0A", x"00", x"18", x"F9", x"F9", x"FF", x"FE", x"F8", x"FB",
	x"00", x"18", x"F8", x"14", x"09", x"EB", x"DA", x"FE", x"F7", x"02", x"10", x"15",
	x"04", x"05", x"0D", x"EF", x"E0", x"01", x"E7", x"F3", x"17", x"16", x"0C", x"16",
	x"05", x"0A", x"EB", x"F3", x"DE", x"E7", x"10", x"03", x"01", x"0C", x"09", x"10",
	x"F7", x"FA", x"F4", x"E9", x"04", x"30", x"17", x"03", x"EC", x"FF", x"EC", x"F3",
	x"C9", x"EA", x"12", x"1A", x"FF", x"11", x"33", x"1C", x"F0", x"EC", x"EE", x"E9",
	x"F5", x"EF", x"28", x"12", x"1D", x"02", x"E2", x"E6", x"DC", x"EF", x"02", x"16",
	x"21", x"F5", x"13", x"0E", x"F2", x"F0", x"FB", x"07", x"FC", x"FD", x"12", x"EF",
	x"0F", x"FF", x"F8", x"F6", x"FF", x"F4", x"00", x"F8", x"16", x"F2", x"27", x"01",
	x"01", x"F0", x"08", x"EE", x"F9", x"E0", x"04", x"01", x"13", x"F2", x"1A", x"FE",
	x"1D", x"F4", x"EE", x"DC", x"23", x"01", x"FE", x"FD", x"16", x"EF", x"F6", x"00",
	x"E9", x"01", x"1F", x"F3", x"05", x"0B", x"F8", x"F5", x"0D", x"FB", x"FF", x"F8",
	x"05", x"E3", x"FF", x"03", x"1A", x"05", x"16", x"F5", x"F6", x"F4", x"EA", x"F8",
	x"FF", x"1A", x"1A", x"01", x"EC", x"12", x"F1", x"08", x"D6", x"06", x"FC", x"06",
	x"03", x"06", x"00", x"13", x"ED", x"F6", x"03", x"F8", x"FF", x"01", x"09", x"28",
	x"10", x"03", x"E1", x"ED", x"D9", x"F3", x"FB", x"1C", x"03", x"2A", x"F4", x"03",
	x"E0", x"0F", x"E7", x"15", x"FE", x"08", x"06", x"03", x"FC", x"ED", x"FD", x"1B",
	x"F5", x"FB", x"F8", x"13", x"ED", x"FD", x"EF", x"FC", x"F9", x"17", x"08", x"0F",
	x"09", x"FD", x"EF", x"F5", x"04", x"FA", x"FC", x"FF", x"14", x"0F", x"EF", x"02",
	x"01", x"DF", x"F7", x"F0", x"04", x"03", x"1C", x"14", x"22", x"0C", x"FC", x"CE",
	x"E9", x"F9", x"EC", x"FF", x"13", x"14", x"0E", x"17", x"00", x"D9", x"EF", x"F5",
	x"F8", x"03", x"2D", x"FE", x"20", x"F0", x"F8", x"CF", x"FA", x"F2", x"1B", x"0D",
	x"09", x"10", x"05", x"ED", x"0C", x"FC", x"ED", x"F2", x"05", x"FD", x"01", x"09",
	x"FF", x"EF", x"25", x"ED", x"ED", x"01", x"07", x"E4", x"0A", x"16", x"08", x"00",
	x"1E", x"03", x"F4", x"EE", x"F1", x"EC", x"10", x"04", x"E7", x"03", x"17", x"FC",
	x"01", x"02", x"F9", x"01", x"04", x"F4", x"00", x"17", x"1D", x"E7", x"07", x"E6",
	x"E4", x"F9", x"00", x"0C", x"10", x"0C", x"03", x"06", x"1D", x"0B", x"E9", x"FD",
	x"E0", x"E7", x"E8", x"FB", x"03", x"0A", x"19", x"05", x"15", x"07", x"F6", x"06",
	x"01", x"F4", x"0B", x"FA", x"F2", x"FA", x"20", x"F0", x"DB", x"FE", x"EB", x"11",
	x"14", x"FB", x"FE", x"25", x"18", x"F5", x"E6", x"F4", x"EE", x"00", x"02", x"E1",
	x"0B", x"1B", x"15", x"0B", x"EC", x"F6", x"04", x"FF", x"DD", x"06", x"14", x"FD",
	x"05", x"0F", x"02", x"1D", x"06", x"EC", x"CB", x"FC", x"FA", x"F6", x"04", x"1A",
	x"08", x"1B", x"EF", x"DC", x"F2", x"07", x"2C", x"F0", x"00", x"FD", x"10", x"10",
	x"F9", x"F7", x"F7", x"04", x"E4", x"F4", x"F7", x"28", x"19", x"02", x"D5", x"00",
	x"FF", x"F8", x"EA", x"05", x"1A", x"08", x"03", x"F5", x"08", x"19", x"10", x"E6",
	x"F2", x"EA", x"03", x"0E", x"0B", x"F5", x"FC", x"01", x"ED", x"EC", x"00", x"2B",
	x"15", x"FD", x"F5", x"FF", x"F5", x"F9", x"F3", x"0D", x"FB", x"F6", x"0B", x"FA",
	x"02", x"14", x"FF", x"EC", x"04", x"05", x"1A", x"F1", x"0E", x"DF", x"FC", x"F6",
	x"F6", x"FF", x"0A", x"1B", x"17", x"E7", x"F1", x"03", x"01", x"05", x"00", x"E1",
	x"05", x"0E", x"0D", x"E8", x"09", x"13", x"08", x"F2", x"F5", x"F8", x"17", x"F4",
	x"FC", x"E8", x"0C", x"01", x"14", x"ED", x"0C", x"FB", x"F9", x"F8", x"05", x"ED",
	x"FF", x"22", x"FC", x"FE", x"07", x"0F", x"FC", x"E7", x"F7", x"F5", x"0D", x"01",
	x"0E", x"08", x"08", x"16", x"FE", x"D4", x"D7", x"09", x"F0", x"04", x"18", x"24",
	x"FB", x"07", x"00", x"ED", x"E3", x"02", x"08", x"F6", x"10", x"13", x"F0", x"0A",
	x"07", x"F6", x"E1", x"00", x"FC", x"0A", x"11", x"2A", x"F2", x"FA", x"DB", x"EC",
	x"F4", x"03", x"02", x"11", x"04", x"1A", x"0A", x"05", x"F1", x"EC", x"EC", x"FE",
	x"05", x"16", x"01", x"11", x"11", x"FB", x"D1", x"E8", x"04", x"01", x"16", x"02",
	x"01", x"F6", x"08", x"01", x"F7", x"FA", x"1B", x"02", x"F5", x"FB", x"04", x"FD",
	x"02", x"01", x"FC", x"E7", x"0F", x"0F", x"EF", x"F2", x"12", x"F8", x"04", x"F0",
	x"F3", x"17", x"24", x"00", x"DF", x"F1", x"15", x"EE", x"F3", x"FB", x"17", x"00",
	x"19", x"06", x"00", x"F0", x"0D", x"D8", x"E1", x"04", x"19", x"14", x"FE", x"11",
	x"00", x"E2", x"FB", x"06", x"F2", x"F8", x"21", x"1B", x"FF", x"F1", x"FA", x"EC",
	x"F0", x"EF", x"EF", x"F4", x"24", x"23", x"0E", x"12", x"0C", x"ED", x"F4", x"EF",
	x"E2", x"FD", x"01", x"07", x"1E", x"0D", x"07", x"F6", x"EA", x"DA", x"DC", x"11",
	x"21", x"16", x"15", x"0B", x"03", x"F2", x"E1", x"D9", x"07", x"12", x"0C", x"06",
	x"0D", x"00", x"02", x"FD", x"01", x"E5", x"EF", x"0B", x"0D", x"F0", x"F5", x"1D",
	x"0C", x"F9", x"FC", x"F4", x"ED", x"0E", x"18", x"E8", x"EC", x"18", x"0E", x"EC",
	x"13", x"08", x"F7", x"FD", x"05", x"EA", x"FB", x"19", x"FA", x"DB", x"07", x"06",
	x"0E", x"0E", x"09", x"EE", x"E8", x"0B", x"04", x"FB", x"12", x"07", x"09", x"F5",
	x"E3", x"F8", x"E3", x"03", x"1A", x"0A", x"13", x"04", x"14", x"F9", x"F2", x"E8",
	x"E2", x"F0", x"20", x"04", x"02", x"1E", x"21", x"E8", x"E4", x"F7", x"F2", x"04",
	x"F8", x"FC", x"0B", x"1B", x"05", x"01", x"F8", x"F0", x"ED", x"F3", x"F4", x"15",
	x"14", x"13", x"20", x"05", x"D3", x"E1", x"F7", x"FF", x"F9", x"06", x"21", x"01",
	x"19", x"F0", x"E4", x"05", x"00", x"02", x"DB", x"14", x"13", x"14", x"00", x"03",
	x"F1", x"09", x"EA", x"ED", x"E7", x"0A", x"1F", x"05", x"11", x"F2", x"06", x"F6",
	x"07", x"05", x"DF", x"F4", x"13", x"04", x"F1", x"0A", x"0B", x"0A", x"03", x"04",
	x"EC", x"03", x"07", x"F6", x"E3", x"FB", x"0D", x"0C", x"19", x"0B", x"EA", x"E6",
	x"01", x"F9", x"0B", x"EC", x"1F", x"15", x"05", x"EF", x"EC", x"FF", x"06", x"00",
	x"F2", x"F4", x"1A", x"0F", x"EE", x"13", x"02", x"EC", x"ED", x"F3", x"EB", x"F7",
	x"41", x"0D", x"05", x"FB", x"0C", x"EC", x"F6", x"E9", x"ED", x"EA", x"38", x"07",
	x"FB", x"07", x"1A", x"19", x"E8", x"D5", x"DB", x"F2", x"17", x"03", x"02", x"26",
	x"0E", x"00", x"F1", x"E8", x"06", x"FA", x"ED", x"FA", x"1D", x"1E", x"09", x"00",
	x"F4", x"DE", x"FC", x"F1", x"FA", x"04", x"11", x"22", x"04", x"04", x"E9", x"EF",
	x"FF", x"F3", x"DE", x"15", x"19", x"17", x"FF", x"0D", x"ED", x"EF", x"F5", x"F6",
	x"03", x"FF", x"13", x"0C", x"FF", x"10", x"FA", x"F8", x"F2", x"0A", x"DD", x"F0",
	x"01", x"21", x"01", x"1A", x"07", x"E9", x"F2", x"FF", x"F1", x"F7", x"0D", x"0B",
	x"02", x"14", x"F9", x"E9", x"01", x"1A", x"FE", x"F4", x"F5", x"10", x"F3", x"EB",
	x"F4", x"0F", x"1A", x"09", x"00", x"FC", x"F1", x"01", x"EC", x"EE", x"F8", x"25",
	x"13", x"FA", x"FE", x"ED", x"07", x"14", x"FE", x"DF", x"06", x"11", x"02", x"FC",
	x"F4", x"03", x"02", x"02", x"E8", x"E6", x"0B", x"32", x"0D", x"F5", x"01", x"04",
	x"EF", x"DE", x"FA", x"EE", x"08", x"16", x"22", x"04", x"06", x"0C", x"F3", x"D9",
	x"EF", x"F0", x"05", x"1B", x"12", x"F5", x"0B", x"17", x"F5", x"D0", x"08", x"07",
	x"01", x"07", x"F5", x"05", x"18", x"FA", x"EE", x"EA", x"FE", x"F3", x"09", x"1B",
	x"0B", x"03", x"0E", x"F0", x"EA", x"E7", x"02", x"00", x"15", x"16", x"F6", x"03",
	x"08", x"02", x"F0", x"F9", x"EF", x"F3", x"07", x"0B", x"0B", x"13", x"F1", x"EF",
	x"FB", x"FA", x"02", x"04", x"FF", x"09", x"F6", x"00", x"FC", x"1F", x"0D", x"00",
	x"FE", x"01", x"D9", x"F5", x"EE", x"02", x"0E", x"1A", x"00", x"F9", x"11", x"02",
	x"E6", x"04", x"ED", x"F4", x"F8", x"11", x"0C", x"04", x"0E", x"11", x"F2", x"FC",
	x"DD", x"03", x"F4", x"09", x"0C", x"0A", x"0F", x"14", x"EC", x"E7", x"EC", x"08",
	x"F6", x"FD", x"1A", x"00", x"08", x"07", x"F7", x"E4", x"FB", x"0C", x"02", x"00",
	x"13", x"F1", x"F9", x"19", x"FD", x"F2", x"FF", x"02", x"EA", x"FC", x"1C", x"F6",
	x"07", x"0D", x"FD", x"FB", x"FF", x"F2", x"FC", x"F2", x"09", x"FC", x"04", x"F5",
	x"00", x"11", x"FC", x"0A", x"09", x"F9", x"F9", x"0D", x"05", x"E9", x"ED", x"16",
	x"FA", x"07", x"07", x"F5", x"FC", x"0B", x"F5", x"E3", x"F8", x"20", x"06", x"FD",
	x"FB", x"00", x"01", x"01", x"00", x"02", x"F2", x"15", x"FC", x"F7", x"FC", x"12",
	x"01", x"F5", x"F9", x"FD", x"E7", x"0F", x"F8", x"F7", x"06", x"1A", x"03", x"FE",
	x"03", x"04", x"F7", x"F7", x"F4", x"02", x"01", x"09", x"FF", x"F8", x"F6", x"05",
	x"04", x"09", x"02", x"0D", x"F3", x"FB", x"FD", x"01", x"04", x"07", x"05", x"ED",
	x"F8", x"01", x"FE", x"F1", x"16", x"08", x"FF", x"F3", x"FC", x"F9", x"04", x"05",
	x"03", x"EB", x"13", x"15", x"FB", x"EE", x"0C", x"03", x"F0", x"01", x"FE", x"02",
	x"09", x"F7", x"EB", x"FD", x"20", x"FB", x"EC", x"03", x"FE", x"F1", x"15", x"F6",
	x"12", x"0B", x"0E", x"E7", x"EC", x"F5", x"FA", x"0F", x"02", x"F9", x"12", x"20",
	x"FA", x"E6", x"EC", x"0C", x"F6", x"F8", x"FD", x"04", x"11", x"13", x"0A", x"F2",
	x"EF", x"FA", x"EA", x"FB", x"12", x"0F", x"FF", x"0D", x"F7", x"FE", x"FD", x"00",
	x"E9", x"F7", x"01", x"15", x"0C", x"0C", x"F8", x"04", x"0F", x"00", x"CB", x"EA",
	x"08", x"21", x"FA", x"F5", x"04", x"12", x"0B", x"FB", x"EF", x"FA", x"FF", x"00",
	x"F4", x"FB", x"12", x"12", x"F9", x"FF", x"05", x"1B", x"ED", x"EF", x"ED", x"F0",
	x"FB", x"03", x"07", x"07", x"10", x"12", x"FD", x"E9", x"09", x"03", x"00", x"06",
	x"FD", x"E4", x"FF", x"1B", x"FA", x"EB", x"06", x"FA", x"00", x"F5", x"0A", x"0B",
	x"1D", x"11", x"F4", x"DC", x"F5", x"E8", x"F7", x"05", x"1D", x"06", x"15", x"14",
	x"FD", x"EB", x"FD", x"E2", x"F0", x"EB", x"19", x"0B", x"0D", x"12", x"15", x"FB",
	x"E8", x"F6", x"EF", x"DF", x"0F", x"10", x"07", x"10", x"17", x"FA", x"EB", x"F1",
	x"FC", x"E5", x"13", x"FA", x"0E", x"16", x"00", x"F7", x"FF", x"07", x"F9", x"EC",
	x"02", x"11", x"FA", x"01", x"F0", x"0A", x"FF", x"FA", x"02", x"F8", x"02", x"0D",
	x"01", x"08", x"EF", x"00", x"F6", x"F8", x"0A", x"F9", x"00", x"0C", x"09", x"06",
	x"FD", x"FB", x"00", x"FC", x"FC", x"EB", x"F1", x"08", x"F7", x"23", x"04", x"05",
	x"F8", x"0B", x"F5", x"FE", x"01", x"F2", x"EA", x"09", x"06", x"04", x"12", x"0F",
	x"FD", x"F3", x"08", x"ED", x"DD", x"FE", x"0B", x"03", x"11", x"19", x"01", x"F2",
	x"02", x"F6", x"ED", x"FA", x"00", x"02", x"15", x"17", x"01", x"ED", x"06", x"02",
	x"E8", x"E2", x"F9", x"0E", x"10", x"04", x"10", x"01", x"08", x"FE", x"E4", x"EF",
	x"0C", x"14", x"F6", x"08", x"0E", x"FC", x"F4", x"FA", x"EA", x"FD", x"F7", x"10",
	x"04", x"00", x"13", x"09", x"00", x"FD", x"F9", x"FC", x"ED", x"FA", x"0A", x"FD",
	x"04", x"14", x"F3", x"FC", x"FB", x"10", x"E2", x"F5", x"00", x"FB", x"04", x"2C",
	x"08", x"FE", x"FB", x"06", x"ED", x"ED", x"FE", x"F3", x"02", x"0D", x"03", x"FC",
	x"FB", x"0C", x"10", x"F1", x"FE", x"0D", x"EF", x"F3", x"0C", x"08", x"EB", x"0C",
	x"1C", x"F2", x"EA", x"05", x"EA", x"F6", x"29", x"0D", x"ED", x"09", x"16", x"DB",
	x"EB", x"01", x"06", x"F8", x"1B", x"FE", x"06", x"07", x"0A", x"E9", x"F9", x"FD",
	x"FE", x"EA", x"03", x"0F", x"16", x"FC", x"FB", x"03", x"00", x"F6", x"06", x"E8",
	x"FD", x"0D", x"07", x"F3", x"1A", x"08", x"E4", x"F2", x"13", x"F2", x"FE", x"05",
	x"16", x"F6", x"FB", x"FE", x"F9", x"F8", x"13", x"02", x"F6", x"F1", x"08", x"0A",
	x"08", x"FD", x"04", x"ED", x"EF", x"08", x"FF", x"02", x"0E", x"13", x"F5", x"ED",
	x"FF", x"FC", x"F2", x"00", x"07", x"06", x"16", x"0D", x"F2", x"F7", x"06", x"F4",
	x"F0", x"F8", x"00", x"11", x"0E", x"0A", x"FA", x"FE", x"E9", x"0A", x"F0", x"F9",
	x"04", x"14", x"05", x"F4", x"F4", x"0B", x"FB", x"13", x"F2", x"F6", x"06", x"0B",
	x"F9", x"EB", x"0F", x"1A", x"F1", x"F3", x"F4", x"F2", x"0C", x"16", x"00", x"00",
	x"06", x"0E", x"DC", x"FC", x"F6", x"00", x"FA", x"12", x"0A", x"0C", x"F7", x"02",
	x"E5", x"FF", x"04", x"0C", x"0A", x"FC", x"F0", x"03", x"07", x"FC", x"FC", x"09",
	x"05", x"FF", x"F7", x"EB", x"00", x"0A", x"04", x"FC", x"FD", x"08", x"05", x"02",
	x"F0", x"09", x"05", x"02", x"F8", x"FB", x"F6", x"05", x"09", x"02", x"F7", x"09",
	x"02", x"E0", x"0E", x"FA", x"08", x"0C", x"FF", x"F0", x"0B", x"0B", x"EA", x"EF",
	x"08", x"12", x"F7", x"00", x"F0", x"01", x"18", x"03", x"F1", x"EF", x"12", x"FA",
	x"05", x"01", x"06", x"01", x"0B", x"EA", x"FA", x"ED", x"F5", x"0D", x"09", x"00",
	x"07", x"17", x"01", x"EE", x"05", x"F8", x"EC", x"F9", x"F2", x"06", x"1A", x"22",
	x"F7", x"FA", x"03", x"F0", x"F4", x"F1", x"FD", x"07", x"17", x"FC", x"F9", x"F4",
	x"11", x"F7", x"FF", x"FE", x"FE", x"08", x"04", x"03", x"F4", x"FF", x"02", x"FB",
	x"F9", x"06", x"00", x"07", x"05", x"F9", x"F5", x"08", x"FD", x"E8", x"04", x"10",
	x"FF", x"FD", x"0F", x"0C", x"0C", x"EA", x"E8", x"DF", x"15", x"16", x"0B", x"03",
	x"FA", x"F0", x"E9", x"05", x"11", x"02", x"03", x"12", x"FE", x"FF", x"E8", x"F8",
	x"FD", x"FD", x"0A", x"F2", x"06", x"18", x"06", x"FC", x"0C", x"EC", x"E6", x"FC",
	x"13", x"FD", x"03", x"0D", x"FC", x"0C", x"03", x"F5", x"DF", x"07", x"F9", x"02",
	x"FC", x"1F", x"05", x"0C", x"E9", x"F9", x"F8", x"FD", x"F1", x"0D", x"0C", x"0A",
	x"FC", x"05", x"FE", x"FA", x"F2", x"FF", x"00", x"02", x"11", x"FF", x"FA", x"01",
	x"F2", x"03", x"F9", x"FD", x"F3", x"15", x"14", x"0D", x"E9", x"F6", x"FE", x"0E",
	x"F7", x"FF", x"FD", x"FF", x"06", x"FF", x"FD", x"FB", x"0E", x"F8", x"FA", x"03",
	x"FA", x"F6", x"04", x"08", x"01", x"F3", x"0D", x"09", x"06", x"FD", x"FC", x"F3",
	x"FA", x"01", x"FA", x"FB", x"14", x"0C", x"FF", x"05", x"02", x"EA", x"F0", x"EB",
	x"06", x"F9", x"19", x"09", x"13", x"03", x"04", x"E9", x"EA", x"F1", x"07", x"03",
	x"12", x"08", x"00", x"01", x"F6", x"02", x"F3", x"F6", x"09", x"FA", x"13", x"04",
	x"00", x"02", x"0A", x"FA", x"E1", x"E9", x"0E", x"01", x"0F", x"0A", x"06", x"F4",
	x"FA", x"F2", x"02", x"05", x"0E", x"F7", x"09", x"00", x"FA", x"04", x"FD", x"FF",
	x"0D", x"F8", x"F7", x"EE", x"FB", x"0C", x"0A", x"03", x"FE", x"F6", x"0C", x"FB",
	x"02", x"F3", x"06", x"FD", x"F8", x"0C", x"08", x"F5", x"01", x"04", x"F8", x"ED",
	x"0A", x"0C", x"FE", x"08", x"09", x"FC", x"F7", x"00", x"FE", x"EE", x"FB", x"0A",
	x"FE", x"08", x"0E", x"F7", x"F8", x"F7", x"02", x"EA", x"04", x"10", x"05", x"14",
	x"0C", x"F0", x"FD", x"00", x"00", x"F3", x"E7", x"05", x"03", x"19", x"08", x"05",
	x"F4", x"F1", x"F3", x"F9", x"F9", x"16", x"12", x"04", x"F1", x"FC", x"04", x"FD",
	x"03", x"FE", x"FF", x"0A", x"05", x"F6", x"ED", x"05", x"13", x"FD", x"F4", x"F9",
	x"F5", x"14", x"06", x"FF", x"F7", x"09", x"02", x"F2", x"F3", x"FF", x"FF", x"0D",
	x"00", x"FF", x"00", x"04", x"0D", x"FE", x"02", x"F7", x"F6", x"08", x"F7", x"EB",
	x"00", x"0D", x"0B", x"04", x"05", x"03", x"06", x"F9", x"E1", x"EF", x"07", x"06",
	x"05", x"0E", x"0F", x"00", x"FA", x"F2", x"F5", x"09", x"00", x"FC", x"06", x"00",
	x"03", x"F6", x"0A", x"08", x"FA", x"F4", x"FD", x"06", x"02", x"F1", x"FD", x"FD",
	x"0C", x"00", x"F5", x"06", x"07", x"03", x"FB", x"F6", x"06", x"05", x"06", x"00",
	x"F8", x"F3", x"FD", x"10", x"05", x"FC", x"00", x"03", x"FE", x"EC", x"F2", x"01",
	x"18", x"14", x"F9", x"E5", x"F9", x"07", x"02", x"F9", x"0F", x"09", x"05", x"F7",
	x"F2", x"F7", x"04", x"05", x"04", x"FA", x"FB", x"01", x"0C", x"04", x"EB", x"FD",
	x"12", x"08", x"F8", x"F6", x"FC", x"10", x"00", x"EA", x"F6", x"0C", x"13", x"EF",
	x"F1", x"F8", x"0F", x"12", x"07", x"FD", x"00", x"0D", x"F6", x"F0", x"F2", x"F8",
	x"08", x"0D", x"FD", x"FD", x"F1", x"FE", x"0D", x"00", x"00", x"02", x"0B", x"FE",
	x"F3", x"03", x"07", x"FF", x"04", x"EB", x"EE", x"0B", x"11", x"05", x"F7", x"02",
	x"FC", x"0A", x"02", x"F3", x"F5", x"09", x"09", x"F8", x"F2", x"01", x"07", x"03",
	x"FA", x"04", x"FA", x"08", x"0F", x"FD", x"F5", x"FD", x"FF", x"02", x"F0", x"FC",
	x"05", x"0F", x"06", x"F6", x"F8", x"06", x"FF", x"09", x"FA", x"FC", x"FB", x"05",
	x"01", x"F4", x"FA", x"04", x"06", x"FB", x"F4", x"06", x"19", x"06", x"F9", x"EF",
	x"FD", x"0C", x"FF", x"02", x"F6", x"01", x"07", x"03", x"FA", x"02", x"FB", x"FC",
	x"F4", x"FE", x"F1", x"09", x"18", x"07", x"FC", x"EF", x"FA", x"FA", x"02", x"08",
	x"16", x"04", x"03", x"EF", x"F4", x"F1", x"06", x"00", x"03", x"01", x"08", x"03",
	x"01", x"04", x"FE", x"F2", x"F4", x"05", x"F7", x"FA", x"06", x"07", x"09", x"05",
	x"0D", x"EF", x"05", x"F9", x"F3", x"F9", x"0F", x"FC", x"F9", x"0A", x"0A", x"E9",
	x"FB", x"05", x"09", x"04", x"05", x"F9", x"03", x"04", x"FE", x"E9", x"06", x"03",
	x"F5", x"FA", x"FE", x"0A", x"11", x"02", x"FA", x"FE", x"02", x"F9", x"F7", x"05",
	x"04", x"01", x"0C", x"F7", x"01", x"01", x"F8", x"0C", x"FA", x"EC", x"EB", x"14",
	x"06", x"F1", x"00", x"0F", x"09", x"08", x"F3", x"ED", x"09", x"0C", x"FC", x"04",
	x"0C", x"05", x"F5", x"FD", x"EB", x"F2", x"01", x"06", x"F4", x"0C", x"11", x"10",
	x"04", x"FA", x"E6", x"F4", x"0F", x"01", x"EC", x"08", x"08", x"0F", x"FF", x"F9",
	x"F3", x"07", x"0B", x"EF", x"F8", x"0D", x"09", x"F4", x"FD", x"06", x"00", x"0A",
	x"FD", x"F4", x"ED", x"06", x"09", x"03", x"03", x"0F", x"05", x"F5", x"F0", x"EE",
	x"F6", x"0B", x"13", x"FA", x"FC", x"0F", x"0B", x"FA", x"F4", x"FC", x"06", x"02",
	x"F6", x"ED", x"FC", x"19", x"13", x"FC", x"FB", x"FF", x"FA", x"EF", x"F4", x"01",
	x"02", x"0E", x"06", x"08", x"04", x"FA", x"FD", x"F1", x"F1", x"03", x"08", x"09",
	x"02", x"01", x"03", x"07", x"01", x"ED", x"EC", x"05", x"02", x"FF", x"FC", x"08",
	x"13", x"0C", x"FE", x"F6", x"EE", x"F8", x"F9", x"04", x"06", x"07", x"0B", x"FC",
	x"F8", x"F9", x"FA", x"FC", x"10", x"07", x"02", x"FF", x"FE", x"F2", x"F2", x"00",
	x"06", x"F8", x"12", x"09", x"F8", x"FC", x"04", x"FB", x"0A", x"0E", x"F4", x"E6",
	x"03", x"F9", x"F4", x"09", x"05", x"06", x"08", x"0C", x"03", x"F3", x"FA", x"FA",
	x"00", x"F7", x"02", x"F7", x"08", x"FE", x"0B", x"F9", x"06", x"FE", x"05", x"FF",
	x"0E", x"FB", x"ED", x"F6", x"07", x"01", x"FD", x"08", x"FE", x"F4", x"03", x"FF",
	x"F9", x"0A", x"15", x"FA", x"EC", x"FC", x"FD", x"FB", x"0C", x"04", x"05", x"08",
	x"FC", x"EE", x"00", x"F6", x"00", x"FB", x"0E", x"04", x"FF", x"08", x"FB", x"F5",
	x"F8", x"FC", x"0F", x"0E", x"01", x"FA", x"FF", x"F4", x"F7", x"00", x"0A", x"F9",
	x"FF", x"F9", x"F7", x"0F", x"0C", x"00", x"FE", x"06", x"FF", x"E6", x"FF", x"07",
	x"02", x"04", x"FF", x"05", x"F8", x"F9", x"F6", x"0A", x"0A", x"0B", x"F3", x"01",
	x"01", x"01", x"F5", x"F8", x"04", x"F7", x"08", x"09", x"0D", x"FA", x"FC", x"00",
	x"FF", x"F2", x"F3", x"00", x"0F", x"07", x"FB", x"EF", x"01", x"0E", x"02", x"07",
	x"F5", x"0A", x"FC", x"FD", x"FE", x"08", x"FE", x"08", x"EB", x"EA", x"06", x"0A",
	x"08", x"FE", x"0E", x"04", x"F7", x"F3", x"FE", x"FA", x"03", x"0C", x"FA", x"FB",
	x"FC", x"08", x"04", x"04", x"F3", x"FF", x"0A", x"00", x"00", x"F4", x"02", x"0A",
	x"F9", x"F7", x"FF", x"05", x"FF", x"01", x"01", x"F6", x"06", x"0A", x"0C", x"F6",
	x"01", x"F1", x"F3", x"F8", x"07", x"06", x"09", x"07", x"FD", x"F8", x"FC", x"0A",
	x"02", x"FF", x"F9", x"FD", x"FA", x"02", x"07", x"F0", x"0C", x"00", x"00", x"FC",
	x"05", x"F4", x"01", x"04", x"09", x"F4", x"04", x"00", x"05", x"02", x"F6", x"FA",
	x"05", x"0B", x"01", x"FC", x"FF", x"F9", x"FA", x"F9", x"E9", x"03", x"16", x"01",
	x"FA", x"FF", x"01", x"08", x"0C", x"02", x"00", x"07", x"FD", x"E6", x"F5", x"FF",
	x"06", x"06", x"04", x"F7", x"FF", x"0D", x"FD", x"07", x"FB", x"03", x"FF", x"FA",
	x"ED", x"FE", x"02", x"04", x"08", x"FF", x"FD", x"02", x"11", x"01", x"F0", x"F7",
	x"03", x"01", x"FD", x"01", x"FA", x"04", x"0C", x"04", x"F9", x"09", x"07", x"F6",
	x"F4", x"FF", x"FC", x"F6", x"01", x"0B", x"F4", x"06", x"03", x"00", x"FB", x"02",
	x"FD", x"02", x"0B", x"FB", x"F1", x"F8", x"13", x"02", x"05", x"FB", x"04", x"FA",
	x"02", x"FD", x"FE", x"FE", x"04", x"FC", x"FA", x"F2", x"04", x"05", x"01", x"F9",
	x"FE", x"03", x"0E", x"0A", x"FC", x"F5", x"06", x"06", x"FC", x"F3", x"FD", x"07",
	x"08", x"F3", x"F8", x"FC", x"0B", x"03", x"01", x"F7", x"FD", x"05", x"0A", x"FA",
	x"00", x"01", x"FA", x"FE", x"FE", x"FC", x"FE", x"08", x"00", x"FC", x"01", x"04",
	x"05", x"FC", x"01", x"F4", x"00", x"06", x"00", x"ED", x"0B", x"11", x"FB", x"E9",
	x"FB", x"0E", x"03", x"0C", x"F4", x"EB", x"F7", x"0D", x"02", x"04", x"0B", x"FF",
	x"F9", x"0C", x"01", x"FB", x"F9", x"03", x"00", x"F7", x"FB", x"05", x"00", x"05",
	x"01", x"F5", x"FF", x"F0", x"04", x"00", x"06", x"0C", x"05", x"F4", x"00", x"08",
	x"F0", x"02", x"00", x"FF", x"00", x"15", x"FC", x"FB", x"00", x"03", x"F2", x"FB",
	x"05", x"F5", x"FE", x"05", x"09", x"FE", x"03", x"03", x"04", x"F8", x"F9", x"F7",
	x"FB", x"00", x"05", x"02", x"04", x"0B", x"FC", x"F6", x"07", x"06", x"FC", x"08",
	x"04", x"F8", x"EF", x"F9", x"01", x"04", x"07", x"FB", x"FD", x"FE", x"04", x"02",
	x"06", x"06", x"00", x"FC", x"F7", x"ED", x"04", x"0A", x"F9", x"03", x"03", x"FE",
	x"08", x"0B", x"FB", x"F8", x"FD", x"00", x"FC", x"FF", x"00", x"FF", x"0B", x"02",
	x"F3", x"F9", x"FE", x"00", x"FC", x"FB", x"0A", x"07", x"05", x"FD", x"FB", x"03",
	x"01", x"FC", x"F6", x"03", x"0B", x"07", x"FE", x"F3", x"FB", x"06", x"FC", x"FC",
	x"FA", x"FC", x"03", x"03", x"FE", x"06", x"09", x"04", x"FA", x"F8", x"FD", x"F7",
	x"01", x"08", x"FE", x"00", x"05", x"F7", x"FF", x"03", x"06", x"FD", x"F9", x"F9",
	x"F8", x"12", x"07", x"F8", x"F8", x"02", x"FF", x"F8", x"F8", x"FA", x"08", x"14",
	x"04", x"F8", x"06", x"FB", x"FD", x"FC", x"F9", x"FF", x"10", x"F8", x"F7", x"0C",
	x"0C", x"F4", x"04", x"F5", x"F6", x"F5", x"08", x"F9", x"05", x"0A", x"0A", x"FB",
	x"05", x"F3", x"F9", x"08", x"00", x"F5", x"00", x"06", x"04", x"FF", x"03", x"F8",
	x"0F", x"F7", x"FB", x"F9", x"04", x"03", x"03", x"F8", x"00", x"FE", x"09", x"00",
	x"F2", x"00", x"00", x"F7", x"00", x"08", x"0C", x"F8", x"0B", x"05", x"F7", x"F6",
	x"FC", x"08", x"03", x"04", x"FD", x"F5", x"FC", x"06", x"F7", x"04", x"00", x"F7",
	x"FE", x"05", x"0F", x"FF", x"FE", x"FD", x"EF", x"03", x"FE", x"0F", x"01", x"04",
	x"FE", x"01", x"F5", x"01", x"F6", x"FF", x"00", x"05", x"F7", x"FB", x"0A", x"0F",
	x"FB", x"02", x"F4", x"03", x"0C", x"00", x"F1", x"FE", x"FF", x"03", x"FE", x"FF",
	x"00", x"FF", x"00", x"05", x"F9", x"01", x"FC", x"0F", x"06", x"FD", x"FB", x"02",
	x"F3", x"FE", x"FC", x"00", x"01", x"02", x"FE", x"FD", x"0E", x"FC", x"F9", x"F9",
	x"03", x"FC", x"03", x"05", x"08", x"01", x"01", x"FC", x"F1", x"00", x"FE", x"05",
	x"FA", x"FF", x"08", x"02", x"F9", x"09", x"0C", x"EC", x"FD", x"FA", x"F7", x"05",
	x"16", x"F6", x"FF", x"07", x"F9", x"F0", x"FE", x"02", x"06", x"0A", x"08", x"F9",
	x"FF", x"FD", x"FB", x"EE", x"02", x"0A", x"09", x"FB", x"F0", x"0B", x"06", x"01",
	x"02", x"FA", x"FA", x"10", x"05", x"EA", x"F5", x"03", x"0B", x"FC", x"05", x"F1",
	x"FC", x"08", x"06", x"F6", x"FE", x"13", x"07", x"F9", x"FE", x"FC", x"00", x"FF",
	x"FD", x"F7", x"FA", x"04", x"0B", x"F7", x"04", x"11", x"FB", x"F4", x"F7", x"F8",
	x"FF", x"05", x"05", x"F3", x"0C", x"0F", x"09", x"F7", x"FB", x"EF", x"02", x"02",
	x"03", x"FF", x"04", x"0A", x"FE", x"F9", x"EF", x"FC", x"02", x"F9", x"03", x"12",
	x"08", x"FC", x"0A", x"F1", x"F8", x"FA", x"00", x"FA", x"09", x"06", x"FF", x"06",
	x"07", x"F0", x"FD", x"FC", x"01", x"F8", x"00", x"04", x"0A", x"05", x"FF", x"FF",
	x"FD", x"FA", x"FB", x"FF", x"F4", x"10", x"04", x"FB", x"FE", x"04", x"FA", x"F7",
	x"07", x"02", x"F8", x"02", x"06", x"FD", x"05", x"FF", x"02", x"FE", x"05", x"F6",
	x"F6", x"03", x"00", x"FE", x"FB", x"03", x"02", x"03", x"FD", x"01", x"F9", x"FA",
	x"08", x"09", x"FF", x"04", x"FD", x"F5", x"FE", x"0A", x"F6", x"FE", x"06", x"03",
	x"F7", x"05", x"FC", x"04", x"08", x"FD", x"F6", x"FC", x"01", x"FC", x"FE", x"FA",
	x"05", x"06", x"04", x"07", x"FE", x"01", x"F6", x"FA", x"F8", x"02", x"11", x"07",
	x"FE", x"F7", x"FB", x"05", x"02", x"F8", x"F1", x"FD", x"09", x"05", x"F7", x"09",
	x"03", x"0D", x"F8", x"F8", x"F2", x"FF", x"02", x"09", x"FF", x"00", x"03", x"FE",
	x"FD", x"FB", x"09", x"FD", x"F6", x"02", x"FF", x"08", x"05", x"02", x"FB", x"F8",
	x"F5", x"F9", x"01", x"05", x"03", x"0D", x"08", x"F2", x"FB", x"FE", x"05", x"01",
	x"F0", x"FD", x"0A", x"04", x"FC", x"07", x"02", x"FA", x"FE", x"FD", x"FE", x"FE",
	x"0D", x"FE", x"FF", x"FC", x"FF", x"F3", x"FF", x"04", x"FE", x"01", x"FE", x"F7",
	x"07", x"05", x"04", x"FF", x"01", x"FA", x"04", x"FB", x"04", x"FB", x"05", x"F4",
	x"FC", x"00", x"05", x"03", x"0D", x"F1", x"F5", x"02", x"0B", x"FD", x"01", x"02",
	x"F9", x"FF", x"07", x"F8", x"FE", x"04", x"06", x"F3", x"F9", x"0B", x"08", x"07",
	x"06", x"F9", x"F1", x"FC", x"FC", x"F7", x"03", x"0E", x"FF", x"FD", x"07", x"FD",
	x"05", x"FE", x"F7", x"F4", x"FD", x"0E", x"02", x"09", x"F7", x"01", x"02", x"FB",
	x"F0", x"04", x"06", x"09", x"01", x"FF", x"F2", x"07", x"0A", x"FA", x"F8", x"08",
	x"F9", x"04", x"FB", x"03", x"FB", x"03", x"FB", x"F8", x"FF", x"05", x"02", x"08",
	x"02", x"FE", x"00", x"F8", x"FF", x"08", x"FD", x"FD", x"FF", x"FF", x"EE", x"0A",
	x"06", x"FE", x"FD", x"06", x"FA", x"03", x"0E", x"FA", x"F6", x"00", x"F9", x"F6",
	x"0A", x"04", x"02", x"0B", x"05", x"FB", x"F3", x"FC", x"F8", x"FC", x"01", x"04",
	x"0B", x"04", x"02", x"F8", x"FC", x"F6", x"FE", x"03", x"FE", x"0B", x"06", x"09",
	x"F5", x"FB", x"F7", x"FC", x"01", x"FD", x"01", x"02", x"04", x"FF", x"06", x"F8",
	x"05", x"FA", x"00", x"03", x"FC", x"04", x"FB", x"09", x"FF", x"FF", x"FE", x"FB",
	x"F7", x"03", x"00", x"FC", x"07", x"03", x"FB", x"04", x"06", x"F5", x"FA", x"05",
	x"FF", x"05", x"01", x"FE", x"04", x"06", x"FA", x"F6", x"FF", x"FF", x"FF", x"FC",
	x"05", x"FF", x"03", x"FB", x"FE", x"09", x"07", x"02", x"F5", x"00", x"FD", x"FE",
	x"FE", x"FD", x"05", x"00", x"06", x"F7", x"00", x"F9", x"06", x"F9", x"01", x"02",
	x"FC", x"03", x"0B", x"FF", x"F7", x"06", x"00", x"F7", x"FB", x"06", x"FF", x"00",
	x"06", x"F4", x"02", x"05", x"04", x"EC", x"01", x"04", x"04", x"01", x"04", x"02",
	x"09", x"F8", x"F9", x"F9", x"04", x"FD", x"02", x"FE", x"05", x"00", x"04", x"FB",
	x"FA", x"FA", x"FB", x"04", x"FC", x"FC", x"08", x"11", x"06", x"F9", x"FC", x"FA",
	x"01", x"FC", x"FD", x"F4", x"0C", x"04", x"03", x"FB", x"05", x"02", x"FD", x"FC",
	x"EF", x"03", x"02", x"04", x"07", x"03", x"02", x"FF", x"F6", x"FB", x"02", x"01",
	x"FA", x"FE", x"02", x"05", x"0A", x"01", x"F8", x"F8", x"FD", x"01", x"00", x"00",
	x"01", x"07", x"0C", x"FD", x"F8", x"F9", x"FE", x"01", x"F5", x"01", x"FB", x"0A",
	x"05", x"0D", x"F6", x"00", x"F4", x"01", x"F5", x"04", x"08", x"FF", x"02", x"05",
	x"03", x"01", x"07", x"F3", x"FC", x"FE", x"FE", x"F2", x"FE", x"0B", x"00", x"07",
	x"FD", x"FE", x"FB", x"07", x"FC", x"FD", x"03", x"00", x"FF", x"05", x"01", x"01",
	x"FF", x"FA", x"FA", x"F6", x"00", x"0A", x"05", x"02", x"03", x"F8", x"00", x"FE",
	x"F9", x"FB", x"05", x"FE", x"01", x"FF", x"0B", x"03", x"FB", x"F9", x"F2", x"03",
	x"04", x"FB", x"0B", x"0B", x"05", x"FA", x"00", x"F6", x"FA", x"00", x"03", x"F2",
	x"FF", x"05", x"0F", x"09", x"FF", x"F6", x"F5", x"FE", x"FD", x"F9", x"FE", x"07",
	x"15", x"02", x"F4", x"FB", x"03", x"FE", x"05", x"FE", x"FB", x"FD", x"08", x"F7",
	x"00", x"09", x"FD", x"F8", x"06", x"FB", x"01", x"00", x"FD", x"F2", x"02", x"0B",
	x"05", x"F9", x"02", x"F8", x"08", x"02", x"FB", x"FA", x"08", x"09", x"02", x"FD",
	x"F1", x"FE", x"0B", x"FA", x"F8", x"FE", x"03", x"0A", x"04", x"FD", x"FD", x"FD",
	x"03", x"F2", x"FA", x"06", x"00", x"07", x"03", x"02", x"FE", x"FF", x"FF", x"F3",
	x"01", x"FF", x"08", x"00", x"FC", x"07", x"06", x"FB", x"FD", x"F7", x"F7", x"08",
	x"FC", x"04", x"F5", x"09", x"04", x"FC", x"FA", x"03", x"01", x"FE", x"FE", x"00",
	x"FE", x"03", x"03", x"04", x"02", x"05", x"FE", x"FA", x"F1", x"03", x"FE", x"02",
	x"06", x"01", x"FA", x"00", x"FC", x"02", x"FD", x"03", x"02", x"FE", x"FD", x"FE",
	x"04", x"02", x"FA", x"00", x"FD", x"02", x"F9", x"FE", x"04", x"08", x"08", x"FB",
	x"F7", x"FE", x"02", x"02", x"FA", x"F8", x"00", x"06", x"01", x"02", x"FC", x"03",
	x"FE", x"FD", x"FA", x"03", x"04", x"FF", x"01", x"F8", x"06", x"FE", x"09", x"F9",
	x"02", x"04", x"FF", x"F2", x"F6", x"02", x"01", x"02", x"06", x"F6", x"01", x"09",
	x"04", x"F8", x"FE", x"FF", x"04", x"FE", x"FE", x"00", x"F9", x"03", x"07", x"F8",
	x"FD", x"01", x"06", x"FB", x"04", x"F6", x"05", x"01", x"07", x"FC", x"FA", x"00",
	x"FA", x"FD", x"06", x"03", x"04", x"04", x"FA", x"F8", x"FA", x"02", x"03", x"FE",
	x"06", x"FE", x"06", x"FE", x"00", x"FC", x"FB", x"FE", x"FF", x"01", x"03", x"00",
	x"07", x"01", x"F8", x"FE", x"F8", x"00", x"02", x"FE", x"FD", x"FE", x"02", x"08",
	x"FB", x"FE", x"04", x"02", x"FD", x"F6", x"03", x"03", x"07", x"05", x"F3", x"F8",
	x"02", x"04", x"FE", x"FE", x"04", x"00", x"03", x"F9", x"F7", x"00", x"01", x"03",
	x"04", x"02", x"00", x"01", x"FD", x"03", x"F8", x"FD", x"00", x"03", x"00", x"FE",
	x"03", x"FC", x"FD", x"FE", x"06", x"01", x"03", x"FE", x"FD", x"04", x"03", x"01",
	x"EF", x"03", x"FD", x"FB", x"02", x"00", x"06", x"08", x"FD", x"FA", x"FD", x"FA",
	x"FF", x"09", x"FE", x"FF", x"FC", x"05", x"FC", x"03", x"00", x"FE", x"F8", x"01",
	x"00", x"02", x"05", x"F8", x"FD", x"06", x"FC", x"FC", x"F9", x"09", x"03", x"0B",
	x"F6", x"FC", x"FC", x"03", x"FE", x"02", x"FF", x"03", x"01", x"00", x"00", x"FF",
	x"00", x"FB", x"F4", x"03", x"FE", x"03", x"02", x"FC", x"04", x"01", x"FF", x"01",
	x"FF", x"FC", x"03", x"06", x"FE", x"F4", x"01", x"FF", x"00", x"01", x"00", x"00",
	x"08", x"00", x"FA", x"FB", x"05", x"00", x"FE", x"00", x"04", x"FA", x"FD", x"F9",
	x"FD", x"FF", x"0C", x"FB", x"00", x"F8", x"07", x"05", x"02", x"FE", x"00", x"FD",
	x"FF", x"F8", x"FD", x"02", x"05", x"FD", x"02", x"FD", x"FE", x"FC", x"05", x"00",
	x"04", x"FA", x"F7", x"F8", x"04", x"06", x"05", x"01", x"FD", x"FF", x"0A", x"FA",
	x"04", x"F8", x"FD", x"FF", x"00", x"FC", x"02", x"05", x"02", x"FE", x"FE", x"02",
	x"FA", x"04", x"F8", x"FD", x"02", x"04", x"02", x"FC", x"05", x"FD", x"FE", x"FC",
	x"F6", x"03", x"07", x"04", x"02", x"FF", x"03", x"FE", x"FB", x"FE", x"F4", x"02",
	x"08", x"04", x"FD", x"03", x"04", x"FE", x"F3", x"F8", x"00", x"05", x"02", x"06",
	x"FF", x"FE", x"01", x"FB", x"FB", x"04", x"FD", x"FB", x"FF", x"04", x"02", x"05",
	x"08", x"01", x"FA", x"FC", x"F2", x"FB", x"04", x"07", x"FD", x"FE", x"04", x"00",
	x"FA", x"02", x"FA", x"FE", x"05", x"FD", x"FF", x"02", x"0B", x"05", x"FD", x"F9",
	x"F7", x"F9", x"02", x"06", x"FB", x"02", x"FF", x"00", x"01", x"05", x"FB", x"00",
	x"00", x"F7", x"FE", x"04", x"0B", x"FA", x"FC", x"00", x"FF", x"FD", x"09", x"F8",
	x"03", x"06", x"05", x"F7", x"FD", x"FE", x"02", x"02", x"FA", x"F7", x"04", x"05",
	x"05", x"FC", x"FC", x"FF", x"FD", x"07", x"02", x"FD", x"FC", x"FF", x"FF", x"F7",
	x"04", x"03", x"06", x"F8", x"08", x"FE", x"F7", x"04", x"05", x"F6", x"04", x"03",
	x"FE", x"FB", x"FE", x"FE", x"FD", x"02", x"FE", x"FB", x"FF", x"06", x"04", x"01",
	x"FF", x"00", x"FD", x"FE", x"FE", x"F9", x"00", x"05", x"00", x"01", x"01", x"01",
	x"03", x"F9", x"00", x"FF", x"FE", x"02", x"FD", x"03", x"FD", x"04", x"F9", x"FA",
	x"FA", x"03", x"04", x"09", x"FD", x"00", x"FC", x"05", x"00", x"FF", x"FE", x"FC",
	x"06", x"FE", x"FD", x"02", x"FE", x"02", x"03", x"FE", x"FA", x"F4", x"FC", x"05",
	x"00", x"06", x"03", x"0B", x"F9", x"05", x"FD", x"F3", x"FB", x"05", x"03", x"03",
	x"FC", x"04", x"FE", x"05", x"FE", x"F6", x"FF", x"02", x"FC", x"00", x"01", x"00",
	x"FE", x"FC", x"05", x"FB", x"06", x"03", x"FC", x"FA", x"07", x"07", x"FA", x"FE",
	x"00", x"01", x"FE", x"FA", x"F9", x"00", x"04", x"0E", x"FA", x"F6", x"04", x"FE",
	x"02", x"01", x"F8", x"FA", x"06", x"07", x"F8", x"FE", x"05", x"00", x"03", x"FE",
	x"FE", x"FE", x"03", x"FC", x"F9", x"FA", x"03", x"02", x"08", x"00", x"04", x"02",
	x"FD", x"F5", x"FA", x"FF", x"04", x"02", x"06", x"FF", x"FF", x"FD", x"01", x"FD",
	x"FE", x"FD", x"FC", x"FB", x"09", x"08", x"05", x"01", x"FA", x"FC", x"F8", x"00",
	x"FD", x"FB", x"04", x"06", x"04", x"FC", x"06", x"FB", x"F9", x"01", x"02", x"F9",
	x"00", x"02", x"0A", x"03", x"00", x"F5", x"F7", x"FD", x"0D", x"04", x"F9", x"FF",
	x"02", x"FF", x"05", x"F9", x"FB", x"FB", x"06", x"04", x"F8", x"00", x"08", x"02",
	x"01", x"FA", x"F9", x"00", x"08", x"01", x"00", x"F8", x"02", x"00", x"FB", x"FD",
	x"04", x"00", x"00", x"FF", x"FC", x"00", x"0B", x"FE", x"F9", x"FE", x"06", x"00",
	x"FD", x"00", x"00", x"F5", x"02", x"FD", x"00", x"03", x"0A", x"05", x"FC", x"FC",
	x"FF", x"FC", x"FD", x"FB", x"03", x"FA", x"04", x"06", x"01", x"FA", x"03", x"01",
	x"FB", x"FB", x"00", x"03", x"03", x"09", x"FC", x"FB", x"FF", x"04", x"FB", x"00",
	x"F7", x"FF", x"04", x"06", x"00", x"FF", x"FF", x"FE", x"FF", x"F9", x"FC", x"08",
	x"02", x"0A", x"01", x"FA", x"F5", x"03", x"FF", x"FB", x"FD", x"0D", x"FD", x"03",
	x"FF", x"01", x"FB", x"04", x"FD", x"F7", x"FA", x"07", x"00", x"01", x"FF", x"0B",
	x"FD", x"FF", x"FC", x"FF", x"01", x"06", x"FA", x"F8", x"F9", x"08", x"07", x"F7",
	x"FE", x"FF", x"00", x"01", x"00", x"FD", x"FE", x"05", x"07", x"FE", x"00", x"FC",
	x"FE", x"FB", x"FE", x"FF", x"FE", x"02", x"06", x"FA", x"FE", x"FF", x"03", x"FC",
	x"03", x"04", x"FF", x"F9", x"06", x"F6", x"04", x"02", x"05", x"F8", x"FE", x"FE",
	x"FD", x"FF", x"03", x"00", x"FE", x"02", x"FF", x"FF", x"FD", x"FD", x"FF", x"FA",
	x"09", x"01", x"01", x"FC", x"05", x"08", x"01", x"F4", x"FE", x"F8", x"FF", x"FE",
	x"FF", x"FD", x"0B", x"04", x"FD", x"FC", x"01", x"02", x"F8", x"F7", x"FE", x"0B",
	x"02", x"05", x"FF", x"02", x"00", x"02", x"F6", x"F4", x"FE", x"0A", x"04", x"00",
	x"FF", x"FE", x"01", x"04", x"F7", x"F6", x"02", x"06", x"06", x"01", x"FE", x"FE",
	x"01", x"01", x"F6", x"F9", x"04", x"07", x"FE", x"04", x"00", x"01", x"00", x"FA",
	x"FA", x"03", x"02", x"00", x"FD", x"FB", x"04", x"03", x"00", x"F8", x"FF", x"05",
	x"FF", x"FB", x"F8", x"01", x"06", x"03", x"FF", x"FA", x"07", x"07", x"FE", x"F7",
	x"FB", x"FC", x"03", x"02", x"04", x"03", x"FF", x"FD", x"FF", x"FB", x"FE", x"FC",
	x"05", x"FF", x"04", x"FD", x"FE", x"FF", x"05", x"FD", x"02", x"FF", x"FE", x"FA",
	x"03", x"04", x"FA", x"02", x"04", x"04", x"03", x"FA", x"FA", x"FB", x"02", x"04",
	x"01", x"01", x"01", x"F9", x"F7", x"FB", x"FE", x"0C", x"03", x"00", x"00", x"02",
	x"FE", x"FC", x"FE", x"FC", x"05", x"02", x"FA", x"04", x"03", x"06", x"04", x"F8",
	x"F9", x"FC", x"FD", x"FC", x"F5", x"04", x"05", x"06", x"FE", x"02", x"FF", x"03",
	x"00", x"FB", x"F8", x"02", x"06", x"07", x"FD", x"FD", x"FD", x"FF", x"FF", x"FD",
	x"FD", x"FE", x"02", x"06", x"01", x"FC", x"F7", x"00", x"FE", x"05", x"03", x"03",
	x"02", x"FE", x"FF", x"FC", x"FE", x"FD", x"00", x"02", x"02", x"03", x"FB", x"FB",
	x"03", x"03", x"06", x"F9", x"FC", x"FE", x"00", x"FD", x"03", x"02", x"03", x"00",
	x"FE", x"FF", x"01", x"00", x"FD", x"01", x"FD", x"FA", x"FB", x"03", x"06", x"02",
	x"04", x"FE", x"FE", x"04", x"04", x"F6", x"FC", x"00", x"02", x"FE", x"01", x"FC",
	x"02", x"00", x"03", x"FA", x"00", x"01", x"02", x"FF", x"F6", x"FE", x"04", x"02",
	x"00", x"08", x"03", x"FF", x"FD", x"00", x"F7", x"FB", x"02", x"FB", x"03", x"FF",
	x"04", x"02", x"00", x"01", x"FE", x"FC", x"00", x"FB", x"FC", x"04", x"00", x"07",
	x"F7", x"00", x"01", x"03", x"01", x"02", x"FD", x"FD", x"00", x"FF", x"F8", x"02",
	x"02", x"FB", x"00", x"03", x"FC", x"01", x"01", x"06", x"FF", x"00", x"FE", x"FA",
	x"03", x"01", x"FA", x"FB", x"FC", x"04", x"05", x"02", x"00", x"FF", x"FC", x"03",
	x"F8", x"FB", x"00", x"08", x"05", x"FF", x"FE", x"FE", x"01", x"FE", x"00", x"FA",
	x"F9", x"03", x"06", x"FF", x"03", x"00", x"FC", x"FC", x"FF", x"FE", x"FF", x"FB",
	x"05", x"04", x"03", x"01", x"04", x"FA", x"FB", x"FB", x"FE", x"FD", x"FF", x"03",
	x"07", x"06", x"FF", x"F6", x"FD", x"03", x"04", x"F7", x"00", x"FC", x"02", x"05",
	x"05", x"FF", x"FF", x"FF", x"FD", x"F9", x"FF", x"09", x"04", x"FF", x"FF", x"FE",
	x"FC", x"FD", x"FE", x"FD", x"01", x"01", x"07", x"FF", x"FE", x"04", x"FA", x"FA",
	x"01", x"FD", x"FB", x"01", x"05", x"03", x"02", x"04", x"00", x"FB", x"FE", x"03",
	x"FA", x"FC", x"FF", x"00", x"FF", x"09", x"FE", x"FA", x"05", x"02", x"FB", x"FB",
	x"FC", x"03", x"FF", x"07", x"04", x"FC", x"01", x"FF", x"FB", x"F9", x"FD", x"04",
	x"FE", x"05", x"07", x"FF", x"FC", x"FB", x"FA", x"FE", x"01", x"07", x"F9", x"FC",
	x"07", x"07", x"02", x"FA", x"FE", x"FE", x"FE", x"F9", x"FE", x"00", x"08", x"05",
	x"FF", x"FB", x"F8", x"FF", x"01", x"01", x"02", x"FD", x"04", x"05", x"00", x"FA",
	x"FE", x"07", x"F9", x"FB", x"FD", x"FD", x"00", x"01", x"06", x"FE", x"FD", x"03",
	x"00", x"FD", x"06", x"FF", x"FE", x"F8", x"04", x"05", x"FE", x"FE", x"FE", x"00",
	x"FF", x"00", x"F9", x"FC", x"00", x"05", x"02", x"00", x"FD", x"01", x"02", x"FD",
	x"FC", x"FC", x"04", x"05", x"03", x"03", x"FE", x"F9", x"FA", x"F7", x"FF", x"00",
	x"02", x"05", x"03", x"05", x"FF", x"02", x"F7", x"FD", x"FB", x"F9", x"FF", x"08",
	x"04", x"08", x"01", x"00", x"F7", x"F9", x"FF", x"FD", x"F9", x"01", x"0B", x"08",
	x"01", x"FB", x"00", x"01", x"FC", x"F9", x"F8", x"FE", x"06", x"0D", x"02", x"FE",
	x"FE", x"F9", x"FA", x"FA", x"FC", x"04", x"05", x"04", x"02", x"FE", x"02", x"FB",
	x"FB", x"FC", x"01", x"06", x"02", x"FE", x"01", x"01", x"01", x"01", x"FC", x"F9",
	x"03", x"FF", x"FE", x"FB", x"00", x"01", x"07", x"01", x"FD", x"FA", x"FE", x"FC",
	x"06", x"FB", x"08", x"05", x"02", x"FF", x"F8", x"F7", x"00", x"FC", x"04", x"FD",
	x"06", x"01", x"FD", x"FE", x"07", x"FF", x"FB", x"FD", x"FF", x"F9", x"01", x"07",
	x"FE", x"00", x"02", x"FC", x"FE", x"01", x"09", x"F9", x"FF", x"FE", x"FF", x"00",
	x"02", x"00", x"04", x"F8", x"FE", x"FF", x"FE", x"FD", x"05", x"00", x"02", x"00",
	x"FF", x"F7", x"00", x"FF", x"03", x"00", x"FD", x"06", x"01", x"04", x"FF", x"F9",
	x"F8", x"FF", x"00", x"03", x"00", x"02", x"06", x"FD", x"01", x"FD", x"FB", x"FA",
	x"01", x"FF", x"00", x"02", x"02", x"02", x"04", x"FF", x"F7", x"FB", x"02", x"01",
	x"01", x"07", x"FE", x"FA", x"FF", x"03", x"00", x"00", x"FF", x"00", x"FC", x"FD",
	x"00", x"00", x"01", x"01", x"03", x"F8", x"FD", x"03", x"00", x"FF", x"FF", x"02",
	x"FD", x"FF", x"03", x"FF", x"01", x"07", x"F9", x"FB", x"FE", x"06", x"FB", x"FD",
	x"02", x"03", x"02", x"00", x"FB", x"F9", x"00", x"03", x"02", x"FA", x"07", x"03",
	x"00", x"FA", x"FE", x"FC", x"FE", x"01", x"03", x"FF", x"FF", x"05", x"00", x"FE",
	x"FF", x"FC", x"FB", x"FE", x"FC", x"01", x"03", x"09", x"FF", x"FA", x"FE", x"02",
	x"02", x"FD", x"04", x"F7", x"01", x"FF", x"02", x"FF", x"04", x"01", x"FF", x"FA",
	x"FD", x"02", x"F8", x"03", x"02", x"07", x"01", x"03", x"FC", x"FC", x"F9", x"01",
	x"FD", x"FC", x"0C", x"07", x"FA", x"00", x"FF", x"F6", x"FC", x"04", x"01", x"FE",
	x"08", x"02", x"FE", x"FD", x"02", x"FD", x"F7", x"02", x"03", x"01", x"FF", x"02",
	x"FD", x"02", x"FB", x"FE", x"F9", x"02", x"04", x"01", x"01", x"04", x"FF", x"FF",
	x"02", x"FD", x"F7", x"FD", x"06", x"FE", x"00", x"00", x"03", x"00", x"FF", x"FA",
	x"FA", x"FE", x"08", x"04", x"FE", x"FF", x"FF", x"01", x"FC", x"FF", x"00", x"FE",
	x"03", x"FE", x"FF", x"FF", x"07", x"FE", x"F7", x"FC", x"FE", x"04", x"06", x"FF",
	x"FE", x"03", x"FD", x"02", x"FC", x"00", x"04", x"00", x"FC", x"F6", x"FF", x"04",
	x"00", x"03", x"02", x"FB", x"00", x"03", x"FD", x"FB", x"03", x"02", x"01", x"FC",
	x"FD", x"FF", x"07", x"03", x"FE", x"F8", x"FF", x"03", x"FA", x"01", x"FE", x"07",
	x"01", x"FF", x"FC", x"FF", x"00", x"02", x"FB", x"FE", x"04", x"02", x"FE", x"02",
	x"02", x"FE", x"FF", x"FD", x"FB", x"FD", x"05", x"00", x"01", x"FC", x"04", x"FF",
	x"00", x"FA", x"FA", x"02", x"05", x"08", x"02", x"FE", x"FC", x"FC", x"FB", x"FD",
	x"00", x"03", x"01", x"05", x"03", x"FD", x"FC", x"FB", x"FD", x"00", x"FE", x"FE",
	x"02", x"05", x"07", x"07", x"FD", x"F7", x"FC", x"FF", x"01", x"02", x"00", x"FF",
	x"FC", x"05", x"F8", x"FE", x"04", x"00", x"FD", x"00", x"00", x"02", x"05", x"FF",
	x"FB", x"00", x"00", x"FD", x"FA", x"FD", x"08", x"06", x"FC", x"FD", x"00", x"02",
	x"FF", x"FE", x"FC", x"F8", x"07", x"07", x"F8", x"FD", x"04", x"02", x"02", x"FF",
	x"FA", x"00", x"00", x"FD", x"F6", x"00", x"08", x"06", x"07", x"F6", x"FA", x"FF",
	x"05", x"FA", x"01", x"00", x"04", x"04", x"04", x"F5", x"FC", x"02", x"FA", x"FB",
	x"00", x"04", x"03", x"06", x"03", x"FB", x"FE", x"FF", x"FB", x"FE", x"01", x"03",
	x"01", x"03", x"FD", x"FD", x"02", x"01", x"01", x"FC", x"01", x"FD", x"FD", x"F8",
	x"04", x"06", x"04", x"FF", x"FD", x"FB", x"FF", x"04", x"FF", x"FF", x"FE", x"03",
	x"FF", x"04", x"FF", x"FD", x"FF", x"06", x"FB", x"F8", x"00", x"02", x"04", x"04",
	x"FF", x"F8", x"FC", x"00", x"03", x"FD", x"01", x"00", x"FF", x"03", x"04", x"FE",
	x"FF", x"FE", x"00", x"FD", x"FA", x"FE", x"03", x"FE", x"03", x"04", x"00", x"FE",
	x"FD", x"FD", x"02", x"FF", x"FD", x"FC", x"00", x"05", x"05", x"FD", x"02", x"FA",
	x"FE", x"FD", x"01", x"FD", x"06", x"01", x"04", x"06", x"FD", x"F6", x"FD", x"00",
	x"FE", x"01", x"01", x"FC", x"05", x"02", x"00", x"F9", x"FF", x"FC", x"FC", x"04",
	x"04", x"FF", x"02", x"01", x"FE", x"FF", x"FF", x"01", x"00", x"00", x"FA", x"FE",
	x"03", x"05", x"01", x"F9", x"FD", x"02", x"FE", x"FF", x"01", x"03", x"FF", x"00",
	x"FE", x"FA", x"FE", x"05", x"04", x"F8", x"00", x"FD", x"01", x"00", x"FF", x"FE",
	x"02", x"05", x"FC", x"01", x"FF", x"04", x"FC", x"F9", x"FA", x"06", x"00", x"02",
	x"02", x"FE", x"FF", x"FB", x"FC", x"FD", x"03", x"04", x"01", x"FB", x"01", x"FC",
	x"02", x"02", x"01", x"00", x"01", x"00", x"FF", x"FA", x"FC", x"02", x"03", x"FF",
	x"FA", x"00", x"01", x"05", x"FD", x"FF", x"00", x"00", x"00", x"FE", x"04", x"FD",
	x"FD", x"FF", x"03", x"FA", x"05", x"00", x"00", x"FB", x"02", x"FF", x"00", x"02",
	x"02", x"02", x"FE", x"FD", x"FC", x"FE", x"00", x"01", x"FF", x"FC", x"FF", x"03",
	x"02", x"FB", x"05", x"FE", x"FE", x"FB", x"03", x"00", x"03", x"FA", x"FF", x"FD",
	x"09", x"02", x"01", x"FC", x"FE", x"F8", x"FE", x"01", x"01", x"03", x"01", x"02",
	x"FC", x"FF", x"00", x"00", x"FD", x"FF", x"FD", x"FE", x"07", x"01", x"FC", x"FC",
	x"06", x"FD", x"00", x"FC", x"01", x"02", x"04", x"FC", x"FB", x"FE", x"01", x"05",
	x"FD", x"FC", x"FE", x"03", x"FE", x"01", x"00", x"04", x"FC", x"04", x"FD", x"FC",
	x"FF", x"00", x"FC", x"03", x"02", x"FE", x"00", x"02", x"FB", x"02", x"03", x"01",
	x"FC", x"03", x"FD", x"FE", x"FD", x"FC", x"FE", x"04", x"04", x"01", x"FC", x"03",
	x"FC", x"02", x"01", x"FF", x"FD", x"04", x"FD", x"FF", x"00", x"02", x"04", x"FB",
	x"FF", x"FD", x"FF", x"01", x"02", x"FD", x"00", x"01", x"00", x"FC", x"FB", x"04",
	x"01", x"FE", x"FE", x"04", x"01", x"02", x"03", x"FB", x"FB", x"FD", x"FC", x"FD",
	x"03", x"05", x"00", x"00", x"02", x"FD", x"01", x"FE", x"FF", x"FC", x"00", x"01",
	x"00", x"00", x"02", x"FE", x"FF", x"FF", x"FA", x"FD", x"06", x"04", x"00", x"FE",
	x"FD", x"01", x"FC", x"FD", x"FD", x"02", x"04", x"02", x"02", x"00", x"00", x"00",
	x"FD", x"F7", x"FD", x"FF", x"01", x"01", x"FD", x"01", x"05", x"03", x"FE", x"FC",
	x"FE", x"03", x"FF", x"FD", x"FD", x"06", x"07", x"FF", x"F6", x"F8", x"FF", x"05",
	x"04", x"02", x"01", x"04", x"FE", x"FA", x"FE", x"FB", x"FC", x"03", x"07", x"FE",
	x"FF", x"00", x"01", x"FB", x"00", x"01", x"FE", x"04", x"FE", x"02", x"01", x"03",
	x"F7", x"FA", x"FC", x"0A", x"01", x"FE", x"01", x"FD", x"FE", x"02", x"03", x"F9",
	x"FE", x"01", x"01", x"FE", x"01", x"FE", x"FD", x"02", x"03", x"FE", x"FF", x"02",
	x"00", x"FE", x"FF", x"01", x"FB", x"01", x"FD", x"05", x"FF", x"01", x"FE", x"04",
	x"FE", x"00", x"FD", x"FB", x"FF", x"FD", x"03", x"01", x"05", x"FF", x"00", x"FC",
	x"04", x"FF", x"FD", x"FE", x"FE", x"FE", x"01", x"FF", x"00", x"03", x"FF", x"02",
	x"FB", x"FD", x"FF", x"FF", x"04", x"02", x"FC", x"FE", x"01", x"00", x"FD", x"FD",
	x"01", x"01", x"04", x"FF", x"04", x"FE", x"00", x"FE", x"FD", x"F8", x"04", x"00",
	x"00", x"00", x"02", x"00", x"FD", x"00", x"FD", x"FD", x"FE", x"07", x"FC", x"FF",
	x"04", x"03", x"00", x"FB", x"FD", x"FA", x"02", x"01", x"04", x"FC", x"04", x"06",
	x"00", x"FC", x"F9", x"FC", x"FE", x"04", x"FF", x"FB", x"01", x"03", x"FF", x"FD",
	x"01", x"FF", x"00", x"01", x"00", x"FB", x"02", x"03", x"FD", x"01", x"FE", x"04",
	x"00", x"FD", x"FE", x"FE", x"01", x"FF", x"FF", x"FE", x"01", x"02", x"01", x"F9",
	x"FC", x"02", x"06", x"00", x"03", x"01", x"FB", x"00", x"FE", x"F8", x"00", x"05",
	x"02", x"00", x"00", x"03", x"FC", x"01", x"FE", x"FC", x"FF", x"06", x"FE", x"FB",
	x"00", x"02", x"00", x"FF", x"FF", x"FD", x"FF", x"01", x"02", x"FF", x"FE", x"03",
	x"02", x"FF", x"FE", x"FB", x"FB", x"01", x"02", x"06", x"FE", x"FF", x"00", x"FF",
	x"FA", x"03", x"FD", x"FF", x"02", x"00", x"FE", x"01", x"01", x"00", x"FD", x"01",
	x"FE", x"FC", x"00", x"01", x"FE", x"04", x"03", x"FE", x"F9", x"FE", x"03", x"04",
	x"00", x"FA", x"FE", x"FD", x"00", x"05", x"FB", x"01", x"01", x"01", x"F9", x"FF",
	x"FE", x"01", x"05", x"01", x"FE", x"FE", x"08", x"FE", x"FC", x"F9", x"FC", x"FE",
	x"00", x"03", x"01", x"07", x"05", x"00", x"F9", x"F9", x"FC", x"00", x"01", x"00",
	x"02", x"00", x"04", x"00", x"00", x"FA", x"FC", x"00", x"FE", x"00", x"03", x"03",
	x"03", x"FF", x"FC", x"F9", x"00", x"00", x"FE", x"00", x"06", x"02", x"FE", x"FE",
	x"FD", x"00", x"FA", x"FC", x"FE", x"01", x"0A", x"02", x"04", x"FC", x"00", x"F9",
	x"FF", x"FB", x"01", x"FF", x"04", x"03", x"FD", x"FD", x"00", x"02", x"01", x"FB",
	x"F9", x"00", x"FF", x"07", x"03", x"FE", x"FE", x"00", x"00", x"FD", x"FE", x"FF",
	x"02", x"FD", x"05", x"FD", x"00", x"FD", x"06", x"FC", x"FF", x"FD", x"00", x"02",
	x"02", x"01", x"FE", x"FB", x"FB", x"02", x"03", x"01", x"FC", x"00", x"00", x"02",
	x"00", x"02", x"FE", x"02", x"FC", x"FF", x"FC", x"00", x"02", x"02", x"04", x"FD",
	x"00", x"F9", x"02", x"00", x"01", x"00", x"FC", x"FB", x"03", x"07", x"01", x"02",
	x"F9", x"FF", x"FB", x"02", x"FC", x"00", x"02", x"07", x"02", x"FD", x"FD", x"FF",
	x"03", x"FF", x"FC", x"FC", x"01", x"01", x"01", x"FC", x"FE", x"01", x"FF", x"FD",
	x"01", x"02", x"05", x"01", x"FD", x"F9", x"FE", x"02", x"01", x"00", x"FB", x"02",
	x"02", x"FE", x"00", x"FE", x"00", x"03", x"FB", x"FD", x"02", x"01", x"03", x"FD",
	x"01", x"FD", x"01", x"FF", x"FE", x"FA", x"01", x"02", x"FC", x"FE", x"00", x"05",
	x"02", x"01", x"FA", x"00", x"FD", x"01", x"00", x"FC", x"FF", x"02", x"01", x"FC",
	x"FD", x"03", x"03", x"01", x"FC", x"FC", x"FE", x"00", x"06", x"FD", x"04", x"FF",
	x"FF", x"01", x"FF", x"FE", x"FD", x"FC", x"00", x"03", x"FE", x"06", x"00", x"01",
	x"FC", x"FF", x"FA", x"FF", x"05", x"04", x"FE", x"FF", x"01", x"FD", x"FE", x"02",
	x"01", x"F9", x"02", x"03", x"FD", x"01", x"01", x"00", x"FE", x"FF", x"FC", x"FB",
	x"04", x"03", x"FC", x"03", x"FE", x"02", x"FD", x"02", x"01", x"FE", x"FD", x"FD",
	x"FE", x"01", x"01", x"04", x"02", x"FC", x"02", x"FD", x"FC", x"02", x"FD", x"FE",
	x"01", x"02", x"FE", x"FF", x"00", x"05", x"FB", x"FF", x"FC", x"01", x"FF", x"05",
	x"FF", x"FE", x"FF", x"00", x"01", x"FB", x"FF", x"02", x"02", x"FC", x"03", x"FC",
	x"FF", x"04", x"00", x"F8", x"FD", x"02", x"01", x"03", x"FF", x"FE", x"FD", x"02",
	x"FE", x"FD", x"05", x"03", x"FD", x"FF", x"FF", x"03", x"00", x"FD", x"02", x"FD",
	x"FF", x"FE", x"01", x"FA", x"05", x"00", x"01", x"F8", x"01", x"04", x"07", x"FF",
	x"FB", x"FA", x"F8", x"08", x"01", x"05", x"00", x"05", x"FC", x"FE", x"FA", x"FB",
	x"01", x"03", x"00", x"FA", x"06", x"03", x"03", x"FB", x"01", x"FC", x"FF", x"01",
	x"00", x"FE", x"FF", x"03", x"FD", x"FE", x"FE", x"02", x"FD", x"03", x"FF", x"FF",
	x"FD", x"04", x"FE", x"02", x"FF", x"FF", x"FC", x"FE", x"FE", x"06", x"03", x"FD",
	x"01", x"FA", x"00", x"FC", x"02", x"FE", x"02", x"01", x"00", x"FF", x"01", x"01",
	x"FE", x"FE", x"FC", x"00", x"FD", x"05", x"FF", x"FF", x"FF", x"FC", x"FC", x"00",
	x"FE", x"05", x"02", x"FF", x"00", x"FC", x"04", x"FC", x"00", x"FA", x"02", x"03",
	x"00", x"F9", x"06", x"00", x"FF", x"FE", x"FF", x"FE", x"FE", x"07", x"FD", x"FF",
	x"FE", x"00", x"FC", x"00", x"FF", x"00", x"01", x"03", x"FC", x"FF", x"02", x"FC",
	x"00", x"FC", x"02", x"FF", x"02", x"FF", x"FF", x"00", x"00", x"FD", x"FF", x"02",
	x"00", x"05", x"F9", x"FE", x"FC", x"01", x"FD", x"02", x"FE", x"02", x"03", x"01",
	x"FE", x"FB", x"01", x"FE", x"05", x"00", x"FE", x"FD", x"03", x"FC", x"FB", x"FE",
	x"02", x"00", x"02", x"01", x"03", x"00", x"FD", x"FC", x"FD", x"FF", x"FD", x"FF",
	x"00", x"05", x"FF", x"00", x"FF", x"FD", x"FC", x"FE", x"01", x"00", x"03", x"FD",
	x"03", x"FF", x"01", x"FB", x"FE", x"FD", x"FF", x"01", x"FF", x"03", x"00", x"FF",
	x"FE", x"FF", x"FC", x"FF", x"01", x"01", x"01", x"02", x"FB", x"FE", x"FD", x"FF",
	x"01", x"01", x"03", x"FF", x"FA", x"00", x"01", x"FF", x"01", x"FF", x"FF", x"00",
	x"FF", x"02", x"FE", x"01", x"FD", x"FD", x"FF", x"02", x"FC", x"01", x"FE", x"01",
	x"00", x"03", x"01", x"00", x"00", x"FE", x"FF", x"FD", x"01", x"00", x"FF", x"FD",
	x"FF", x"FA", x"04", x"01", x"03", x"02", x"01", x"FF", x"FF", x"FC", x"FA", x"00",
	x"03", x"03", x"FE", x"01", x"00", x"FF", x"FE", x"00", x"01", x"FD", x"FF", x"00",
	x"00", x"02", x"00", x"FE", x"FE", x"FE", x"01", x"FD", x"04", x"00", x"01", x"FF",
	x"FE", x"F9", x"FF", x"03", x"01", x"00", x"FD", x"00", x"FD", x"04", x"FF", x"02",
	x"FC", x"01", x"FE", x"FF", x"FC", x"01", x"FF", x"FF", x"01", x"FF", x"02", x"FC",
	x"01", x"01", x"FE", x"FF", x"01", x"FB", x"00", x"06", x"FD", x"01", x"FE", x"FE",
	x"FF", x"FF", x"FE", x"FF", x"01", x"05", x"00", x"00", x"00", x"FC", x"FD", x"00",
	x"FA", x"FD", x"04", x"03", x"02", x"00", x"01", x"FC", x"01", x"FA", x"FF", x"FD",
	x"01", x"FE", x"04", x"01", x"02", x"FF", x"00", x"FE", x"FF", x"02", x"FE", x"FF",
	x"FF", x"00", x"00", x"FC", x"FD", x"FD", x"05", x"00", x"04", x"F9", x"FE", x"03",
	x"03", x"FD", x"FF", x"FE", x"01", x"FE", x"02", x"FA", x"FF", x"03", x"04", x"FE",
	x"01", x"FE", x"00", x"FF", x"00", x"FE", x"FB", x"03", x"FD", x"01", x"01", x"02",
	x"00", x"FC", x"FE", x"FF", x"02", x"00", x"03", x"FA", x"00", x"01", x"03", x"FA",
	x"02", x"01", x"FC", x"FF", x"FE", x"03", x"FF", x"03", x"FE", x"FD", x"FF", x"03",
	x"FD", x"00", x"FD", x"FF", x"01", x"02", x"01", x"FF", x"FF", x"04", x"FF", x"FA",
	x"FD", x"FD", x"03", x"FF", x"02", x"00", x"02", x"00", x"00", x"FE", x"FD", x"00",
	x"FF", x"00", x"00", x"03", x"FD", x"01", x"F8", x"FF", x"FD", x"05", x"01", x"06",
	x"FF", x"FD", x"00", x"FE", x"FC", x"00", x"01", x"01", x"02", x"FF", x"00", x"00",
	x"01", x"00", x"FB", x"01", x"FB", x"FF", x"FD", x"05", x"01", x"02", x"00", x"00",
	x"FD", x"02", x"01", x"FE", x"FF", x"01", x"00", x"FF", x"04", x"FF", x"F8", x"FE",
	x"00", x"FF", x"04", x"02", x"00", x"FD", x"03", x"FD", x"FD", x"FE", x"FE", x"02",
	x"00", x"03", x"F9", x"01", x"01", x"05", x"FE", x"FD", x"FB", x"01", x"04", x"01",
	x"FF", x"FA", x"04", x"FE", x"00", x"FB", x"01", x"01", x"02", x"FD", x"FF", x"01",
	x"01", x"01", x"FD", x"FF", x"FD", x"01", x"00", x"FF", x"FF", x"02", x"00", x"FB",
	x"FD", x"03", x"02", x"04", x"FB", x"FF", x"FE", x"00", x"01", x"FD", x"FF", x"01",
	x"05", x"FD", x"FE", x"01", x"02", x"FD", x"FF", x"FC", x"FB", x"03", x"02", x"03",
	x"FE", x"06", x"FF", x"FE", x"FF", x"FE", x"FF", x"03", x"FF", x"FA", x"00", x"00",
	x"02", x"FD", x"FF", x"FE", x"02", x"02", x"02", x"01", x"FF", x"00", x"FC", x"FA",
	x"FD", x"03", x"05", x"00", x"FF", x"01", x"FC", x"00", x"03", x"00", x"FC", x"FD",
	x"01", x"FF", x"02", x"02", x"00", x"00", x"00", x"FD", x"FC", x"FB", x"00", x"02",
	x"03", x"FE", x"FE", x"00", x"02", x"00", x"02", x"FC", x"01", x"03", x"FE", x"FF",
	x"FF", x"01", x"FA", x"FE", x"FD", x"00", x"03", x"01", x"FE", x"FC", x"00", x"00",
	x"FF", x"01", x"01", x"01", x"02", x"02", x"FC", x"FB", x"FC", x"06", x"FD", x"FF",
	x"00", x"FE", x"00", x"00", x"02", x"FD", x"01", x"02", x"FD", x"FD", x"00", x"01",
	x"FF", x"00", x"FE", x"00", x"FF", x"02", x"01", x"FF", x"00", x"FE", x"00", x"FE",
	x"FF", x"00", x"FF", x"00", x"02", x"FE", x"01", x"06", x"FD", x"FB", x"FE", x"FF",
	x"FE", x"FF", x"01", x"01", x"02", x"01", x"02", x"F8", x"FC", x"00", x"00", x"02",
	x"FF", x"00", x"04", x"02", x"00", x"F9", x"FB", x"04", x"00", x"FC", x"00", x"01",
	x"02", x"03", x"01", x"F9", x"FE", x"FE", x"FE", x"FC", x"01", x"07", x"02", x"FD",
	x"FE", x"FE", x"FE", x"01", x"FF", x"FC", x"FE", x"02", x"04", x"FE", x"FE", x"FE",
	x"02", x"FD", x"00", x"FE", x"FE", x"02", x"01", x"FE", x"FE", x"02", x"FF", x"00",
	x"FD", x"00", x"FE", x"01", x"03", x"00", x"FF", x"FD", x"FE", x"FF", x"00", x"03",
	x"FC", x"01", x"00", x"FE", x"FF", x"FE", x"01", x"FD", x"00", x"FF", x"01", x"FA",
	x"03", x"01", x"01", x"00", x"FD", x"00", x"FD", x"01", x"FE", x"02", x"FE", x"05",
	x"FC", x"FF", x"00", x"02", x"FD", x"FB", x"02", x"02", x"00", x"FF", x"02", x"FE",
	x"04", x"02", x"FC", x"FD", x"FF", x"FD", x"00", x"01", x"FE", x"03", x"01", x"FE",
	x"FB", x"00", x"01", x"02", x"FD", x"FC", x"FD", x"03", x"00", x"00", x"FE", x"FF",
	x"02", x"02", x"FD", x"FC", x"00", x"02", x"01", x"FB", x"01", x"FE", x"02", x"FD",
	x"FE", x"FE", x"02", x"03", x"02", x"FD", x"FC", x"06", x"FE", x"FD", x"F9", x"00",
	x"01", x"03", x"02", x"FD", x"07", x"00", x"FE", x"F6", x"FE", x"FE", x"04", x"02",
	x"00", x"FE", x"03", x"04", x"FD", x"FD", x"FC", x"02", x"03", x"FC", x"FF", x"FF",
	x"FF", x"02", x"00", x"FB", x"FD", x"04", x"FF", x"FB", x"FD", x"06", x"03", x"04",
	x"00", x"F9", x"FE", x"FF", x"01", x"FC", x"03", x"00", x"FD", x"FD", x"FD", x"FF",
	x"00", x"02", x"01", x"01", x"FF", x"01", x"00", x"FF", x"FD", x"FF", x"01", x"FC",
	x"FF", x"00", x"03", x"03", x"FF", x"FD", x"01", x"FE", x"FC", x"FE", x"04", x"FE",
	x"00", x"01", x"FF", x"00", x"01", x"00", x"FC", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"01", x"01", x"FE", x"01", x"02", x"01", x"FE", x"00", x"00", x"FE", x"01",
	x"FF", x"FD", x"FF", x"02", x"FF", x"FD", x"00", x"01", x"02", x"01", x"FD", x"FC",
	x"02", x"03", x"FB", x"FB", x"01", x"03", x"00", x"00", x"03", x"FD", x"04", x"00",
	x"FE", x"F9", x"02", x"00", x"FF", x"00", x"FD", x"02", x"00", x"02", x"F8", x"FE",
	x"03", x"01", x"FF", x"FD", x"FF", x"02", x"01", x"00", x"FC", x"00", x"03", x"01",
	x"FC", x"FE", x"00", x"00", x"FC", x"00", x"FE", x"FE", x"03", x"FD", x"01", x"FE",
	x"01", x"FE", x"FE", x"00", x"00", x"06", x"01", x"FE", x"FA", x"FD", x"FD", x"03",
	x"FC", x"03", x"00", x"03", x"FE", x"FF", x"FF", x"FF", x"00", x"FE", x"FB", x"05",
	x"00", x"01", x"00", x"01", x"FA", x"FE", x"FE", x"FF", x"FE", x"04", x"01", x"02",
	x"00", x"FE", x"FF", x"FB", x"FF", x"FC", x"FD", x"02", x"02", x"00", x"01", x"02",
	x"00", x"FC", x"FB", x"01", x"00", x"02", x"00", x"00", x"FE", x"02", x"FE", x"FE",
	x"00", x"00", x"01", x"01", x"01", x"FC", x"FE", x"01", x"02", x"FD", x"FD", x"FE",
	x"01", x"03", x"01", x"FE", x"FE", x"FC", x"FF", x"00", x"04", x"00", x"01", x"FF",
	x"FB", x"01", x"01", x"FF", x"01", x"01", x"01", x"FD", x"FF", x"FE", x"02", x"00",
	x"01", x"FC", x"FF", x"00", x"01", x"FE", x"01", x"FE", x"FF", x"03", x"FD", x"01",
	x"FF", x"04", x"00", x"FE", x"FA", x"00", x"FF", x"FE", x"01", x"03", x"FD", x"04",
	x"02", x"FD", x"00", x"FC", x"FE", x"FB", x"01", x"04", x"01", x"02", x"FF", x"FC",
	x"00", x"FF", x"01", x"FE", x"FF", x"02", x"FF", x"FE", x"FF", x"00", x"01", x"04",
	x"FE", x"FC", x"FD", x"04", x"FD", x"FF", x"00", x"FE", x"02", x"FE", x"01", x"FD",
	x"01", x"FE", x"00", x"FC", x"03", x"02", x"01", x"FE", x"FF", x"02", x"FC", x"FF",
	x"FD", x"00", x"02", x"01", x"00", x"FD", x"03", x"03", x"FF", x"FD", x"FE", x"FC",
	x"00", x"FF", x"FF", x"00", x"05", x"03", x"FD", x"F8", x"FF", x"02", x"02", x"FF",
	x"FF", x"02", x"01", x"01", x"FE", x"FC", x"FE", x"03", x"FE", x"FF", x"00", x"02",
	x"FF", x"00", x"FF", x"FE", x"02", x"00", x"FF", x"FC", x"01", x"01", x"FE", x"FE",
	x"00", x"04", x"FF", x"FE", x"FB", x"FE", x"04", x"03", x"FC", x"FC", x"00", x"02",
	x"FE", x"00", x"FF", x"00", x"02", x"00", x"FF", x"FE", x"00", x"00", x"01", x"FE",
	x"00", x"FF", x"FD", x"FF", x"FD", x"01", x"02", x"02", x"FD", x"FC", x"FE", x"02",
	x"00", x"FF", x"FE", x"00", x"FF", x"02", x"FE", x"01", x"FF", x"FF", x"FD", x"01",
	x"02", x"FE", x"FF", x"FF", x"02", x"FF", x"01", x"FC", x"FF", x"FE", x"02", x"01",
	x"00", x"00", x"FD", x"01", x"FE", x"02", x"FC", x"FF", x"FF", x"03", x"01", x"00",
	x"01", x"FC", x"FB", x"02", x"01", x"00", x"FF", x"FF", x"00", x"03", x"FF", x"FF",
	x"FD", x"FF", x"00", x"01", x"01", x"FD", x"02", x"00", x"FF", x"FC", x"00", x"FF",
	x"02", x"01", x"FE", x"FD", x"00", x"00", x"02", x"02", x"FF", x"FF", x"03", x"FB",
	x"FF", x"01", x"02", x"01", x"FD", x"FE", x"00", x"01", x"01", x"00", x"FF", x"00",
	x"00", x"00", x"FD", x"FE", x"01", x"01", x"FE", x"FD", x"03", x"FD", x"05", x"FE",
	x"FD", x"01", x"03", x"FE", x"FE", x"FF", x"FE", x"03", x"01", x"FE", x"FE", x"05",
	x"02", x"FF", x"FB", x"FD", x"FE", x"02", x"01", x"00", x"FE", x"02", x"01", x"FD",
	x"FE", x"00", x"01", x"FF", x"FB", x"FF", x"02", x"02", x"01", x"FE", x"FC", x"01",
	x"01", x"FD", x"FF", x"03", x"01", x"00", x"FF", x"FE", x"FE", x"FF", x"02", x"FE",
	x"FF", x"00", x"01", x"FC", x"02", x"FE", x"01", x"00", x"FE", x"FC", x"00", x"01",
	x"05", x"FE", x"FE", x"00", x"00", x"01", x"FE", x"FF", x"FD", x"02", x"00", x"FE",
	x"FF", x"FF", x"01", x"FF", x"00", x"FD", x"FF", x"FF", x"02", x"00", x"00", x"FC",
	x"FE", x"01", x"03", x"03", x"FE", x"FC", x"FC", x"01", x"01", x"01", x"FF", x"FF",
	x"FF", x"03", x"00", x"FF", x"FC", x"01", x"FE", x"01", x"FD", x"FF", x"01", x"02",
	x"01", x"FD", x"FA", x"FF", x"02", x"02", x"FF", x"04", x"FD", x"FF", x"FF", x"00",
	x"FC", x"FE", x"FF", x"01", x"FE", x"04", x"FF", x"FF", x"03", x"FF", x"FE", x"FE",
	x"FD", x"FF", x"00", x"04", x"02", x"FE", x"FD", x"02", x"FE", x"FC", x"FC", x"01",
	x"FF", x"05", x"01", x"FD", x"FF", x"05", x"FE", x"FC", x"FD", x"00", x"FF", x"01",
	x"02", x"FE", x"FF", x"03", x"FF", x"FD", x"FD", x"01", x"00", x"FF", x"FF", x"FF",
	x"05", x"01", x"FF", x"FC", x"FD", x"05", x"FD", x"00", x"FF", x"01", x"FE", x"02",
	x"FA", x"00", x"02", x"04", x"FD", x"FE", x"00", x"FF", x"01", x"FD", x"FD", x"00",
	x"02", x"00", x"FE", x"FF", x"02", x"02", x"00", x"FC", x"F9", x"05", x"01", x"01",
	x"FD", x"FF", x"01", x"00", x"FF", x"FE", x"00", x"01", x"01", x"FF", x"00", x"00",
	x"FE", x"FC", x"01", x"00", x"00", x"FF", x"02", x"01", x"01", x"FF", x"FF", x"FA",
	x"00", x"01", x"03", x"FF", x"03", x"FE", x"02", x"00", x"FB", x"FA", x"03", x"04",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"01", x"01", x"00", x"00", x"FE",
	x"FF", x"00", x"FF", x"FD", x"02", x"00", x"00", x"FF", x"FF", x"FE", x"00", x"02",
	x"FF", x"00", x"02", x"01", x"FD", x"FC", x"FF", x"FF", x"05", x"00", x"FD", x"01",
	x"02", x"00", x"FB", x"FC", x"00", x"01", x"00", x"FF", x"00", x"02", x"01", x"02",
	x"FC", x"FA", x"FF", x"FF", x"FE", x"00", x"02", x"02", x"01", x"01", x"FC", x"FC",
	x"00", x"FE", x"01", x"00", x"02", x"00", x"00", x"FF", x"FD", x"02", x"FD", x"FC",
	x"01", x"00", x"00", x"04", x"FF", x"FF", x"FE", x"FF", x"02", x"FD", x"01", x"FF",
	x"FF", x"00", x"FE", x"FD", x"01", x"03", x"01", x"FF", x"FD", x"FE", x"FE", x"02",
	x"FD", x"FF", x"FE", x"00", x"02", x"FF", x"01", x"FE", x"FD", x"00", x"FE", x"FF",
	x"FF", x"02", x"03", x"00", x"FD", x"FF", x"FC", x"FE", x"FE", x"02", x"00", x"01",
	x"00", x"01", x"00", x"01", x"FD", x"FE", x"FD", x"FF", x"FF", x"03", x"02", x"00",
	x"FE", x"00", x"FE", x"00", x"00", x"00", x"FD", x"00", x"FF", x"00", x"00", x"02",
	x"02", x"00", x"FE", x"FF", x"FE", x"00", x"01", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"02", x"FF", x"02", x"FE", x"00", x"FE", x"FE", x"01", x"02", x"01", x"FE", x"FE",
	x"FE", x"03", x"01", x"FE", x"FE", x"00", x"FE", x"FE", x"FD", x"00", x"01", x"01",
	x"01", x"FD", x"00", x"01", x"FF", x"00", x"FE", x"FC", x"00", x"03", x"FF", x"FF",
	x"01", x"01", x"01", x"00", x"FB", x"FD", x"01", x"01", x"FF", x"FF", x"01", x"01",
	x"00", x"00", x"FC", x"02", x"FE", x"01", x"FC", x"01", x"00", x"FF", x"FF", x"FE",
	x"00", x"01", x"02", x"FF", x"00", x"FE", x"04", x"01", x"FF", x"FC", x"00", x"FE",
	x"FE", x"FE", x"00", x"03", x"03", x"02", x"FD", x"FC", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"01", x"01", x"FF", x"00", x"FF", x"FF", x"FC", x"FE", x"02", x"00",
	x"02", x"FF", x"FF", x"FD", x"03", x"00", x"FE", x"FF", x"02", x"00", x"FD", x"FE",
	x"01", x"02", x"FE", x"FF", x"FC", x"00", x"02", x"00", x"01", x"FC", x"FF", x"00",
	x"FE", x"01", x"FE", x"01", x"00", x"FE", x"FF", x"01", x"03", x"FE", x"FF", x"FE",
	x"FE", x"FD", x"04", x"00", x"01", x"02", x"01", x"FD", x"FE", x"00", x"FD", x"00",
	x"FE", x"01", x"00", x"03", x"00", x"01", x"FE", x"FE", x"FC", x"FD", x"FD", x"04",
	x"04", x"00", x"FE", x"FF", x"FE", x"FE", x"03", x"FF", x"00", x"03", x"02", x"FC",
	x"FE", x"00", x"00", x"FF", x"FC", x"FF", x"01", x"03", x"FF", x"FF", x"01", x"00",
	x"FC", x"FD", x"FD", x"03", x"04", x"00", x"FE", x"FE", x"FE", x"04", x"01", x"FD",
	x"FF", x"04", x"00", x"FD", x"01", x"FD", x"00", x"01", x"FE", x"FE", x"FF", x"06",
	x"01", x"FE", x"FB", x"FD", x"02", x"00", x"00", x"00", x"02", x"FF", x"01", x"FE",
	x"00", x"FF", x"01", x"FA", x"FE", x"01", x"01", x"04", x"00", x"01", x"FD", x"FF",
	x"FE", x"FC", x"FD", x"05", x"03", x"00", x"FF", x"FF", x"FE", x"01", x"FF", x"FE",
	x"FF", x"02", x"FF", x"00", x"00", x"01", x"01", x"FC", x"00", x"FE", x"01", x"01",
	x"00", x"00", x"01", x"01", x"FD", x"01", x"FF", x"01", x"FE", x"00", x"FE", x"01",
	x"FE", x"01", x"02", x"FD", x"FF", x"FD", x"FF", x"00", x"FF", x"03", x"02", x"FF",
	x"FF", x"FE", x"00", x"01", x"FE", x"FF", x"00", x"FF", x"FE", x"01", x"FE", x"00",
	x"01", x"FF", x"00", x"FE", x"00", x"01", x"01", x"FD", x"FF", x"FE", x"01", x"FE",
	x"02", x"FE", x"FF", x"FF", x"01", x"FF", x"01", x"FF", x"FE", x"FC", x"01", x"00",
	x"00", x"02", x"FE", x"01", x"00", x"00", x"FC", x"FE", x"FF", x"03", x"00", x"00",
	x"FD", x"02", x"FE", x"01", x"02", x"FC", x"FF", x"FE", x"02", x"FD", x"FF", x"02",
	x"02", x"00", x"FF", x"FC", x"FF", x"02", x"FE", x"02", x"FE", x"00", x"FC", x"00",
	x"FF", x"02", x"00", x"00", x"FE", x"00", x"FE", x"03", x"FE", x"FD", x"FE", x"01",
	x"01", x"01", x"FF", x"01", x"FD", x"FF", x"00", x"FD", x"01", x"FE", x"04", x"FF",
	x"FF", x"02", x"FF", x"FF", x"FD", x"02", x"FF", x"00", x"FF", x"00", x"FE", x"02",
	x"FF", x"FF", x"FC", x"02", x"FF", x"FE", x"02", x"00", x"03", x"01", x"FE", x"FD",
	x"FC", x"FE", x"02", x"FE", x"02", x"00", x"04", x"00", x"FF", x"FC", x"FE", x"FF",
	x"FE", x"FD", x"02", x"03", x"FE", x"00", x"00", x"01", x"FD", x"00", x"FD", x"FF",
	x"01", x"01", x"00", x"FF", x"02", x"00", x"00", x"FC", x"00", x"FE", x"01", x"FE",
	x"02", x"FD", x"02", x"02", x"FF", x"FC", x"FE", x"01", x"00", x"FE", x"FE", x"FF",
	x"01", x"01", x"FB", x"01", x"02", x"01", x"FF", x"FF", x"FD", x"FD", x"02", x"FE",
	x"FE", x"00", x"00", x"FE", x"02", x"FE", x"00", x"01", x"02", x"FD", x"FD", x"00",
	x"FF", x"02", x"FE", x"FF", x"FF", x"03", x"FF", x"01", x"FF", x"00", x"FD", x"FF",
	x"FF", x"01", x"04", x"FE", x"00", x"FD", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"FC", x"03", x"00", x"FF", x"FE", x"02", x"01", x"FF",
	x"FE", x"00", x"FC", x"00", x"FF", x"02", x"02", x"00", x"FE", x"00", x"FF", x"00",
	x"FF", x"FE", x"00", x"01", x"03", x"FF", x"FF", x"FE", x"00", x"01", x"FF", x"00",
	x"FC", x"01", x"01", x"00", x"FC", x"00", x"FD", x"01", x"00", x"02", x"03", x"FF",
	x"01", x"F9", x"FF", x"FE", x"01", x"00", x"FE", x"FF", x"01", x"00", x"FF", x"02",
	x"FF", x"FF", x"FC", x"01", x"FD", x"04", x"02", x"00", x"FE", x"00", x"FE", x"FE",
	x"FE", x"FF", x"00", x"02", x"01", x"FD", x"FF", x"02", x"00", x"FA", x"FD", x"FF",
	x"02", x"04", x"02", x"FF", x"FE", x"00", x"FD", x"FC", x"FA", x"FF", x"03", x"04",
	x"FE", x"03", x"00", x"00", x"FE", x"FC", x"FB", x"FF", x"00", x"FE", x"01", x"01",
	x"02", x"FF", x"03", x"FB", x"00", x"01", x"00", x"FB", x"01", x"02", x"01", x"FF",
	x"FF", x"FD", x"02", x"01", x"FD", x"FF", x"FF", x"02", x"00", x"FD", x"FD", x"01",
	x"02", x"FF", x"01", x"00", x"00", x"FD", x"00", x"FC", x"00", x"FF", x"04", x"FC",
	x"01", x"00", x"FE", x"FF", x"FE", x"FF", x"01", x"00", x"FF", x"FF", x"FF", x"02",
	x"FF", x"FE", x"FD", x"FE", x"01", x"02", x"01", x"FE", x"FF", x"FF", x"FD", x"FE",
	x"FF", x"01", x"02", x"FF", x"01", x"FE", x"00", x"FF", x"FF", x"FE", x"FD", x"01",
	x"02", x"FE", x"00", x"01", x"00", x"FF", x"FC", x"02", x"FB", x"01", x"01", x"FF",
	x"FE", x"00", x"FE", x"01", x"FF", x"FF", x"00", x"FD", x"01", x"01", x"00", x"00",
	x"01", x"FE", x"01", x"FC", x"FD", x"FF", x"00", x"02", x"00", x"01", x"FE", x"FF",
	x"FF", x"03", x"FE", x"FC", x"01", x"FF", x"01", x"02", x"00", x"00", x"FE", x"FF",
	x"FE", x"FD", x"FF", x"00", x"01", x"02", x"01", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"FD", x"02", x"01", x"00", x"02", x"FE", x"00", x"FC", x"01", x"FE", x"01",
	x"FF", x"01", x"00", x"01", x"00", x"FE", x"00", x"FE", x"00", x"00", x"FD", x"02",
	x"01", x"01", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"FC", x"03", x"FF", x"01",
	x"00", x"00", x"FD", x"03", x"FE", x"FF", x"FD", x"01", x"01", x"FF", x"FE", x"02",
	x"FF", x"FF", x"FF", x"FC", x"00", x"00", x"FF", x"FE", x"00", x"02", x"FF", x"FD",
	x"FF", x"FE", x"FE", x"00", x"FF", x"FD", x"00", x"02", x"00", x"00", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"00", x"01", x"FF", x"FF", x"00", x"01", x"03", x"FE",
	x"FF", x"FD", x"00", x"01", x"00", x"00", x"00", x"00", x"FF", x"FE", x"00", x"FE",
	x"02", x"01", x"FE", x"01", x"FF", x"FF", x"FE", x"00", x"01", x"FF", x"FF", x"FF",
	x"FE", x"03", x"02", x"FF", x"FF", x"FC", x"01", x"FF", x"00", x"00", x"FF", x"00",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"01", x"00", x"03", x"FD", x"00", x"00", x"02",
	x"FE", x"FF", x"00", x"FD", x"01", x"01", x"02", x"FE", x"FE", x"FD", x"FF", x"FF",
	x"01", x"FF", x"FF", x"02", x"FF", x"01", x"FF", x"FE", x"00", x"01", x"00", x"FF",
	x"FE", x"01", x"FC", x"02", x"FE", x"00", x"FE", x"00", x"01", x"00", x"01", x"FE",
	x"FF", x"FD", x"00", x"FF", x"03", x"FE", x"02", x"FD", x"04", x"FD", x"FD", x"01",
	x"00", x"02", x"00", x"02", x"FE", x"FF", x"FF", x"FF", x"FB", x"00", x"00", x"00",
	x"02", x"02", x"00", x"FD", x"00", x"FC", x"00", x"FE", x"00", x"FF", x"02", x"01",
	x"00", x"FE", x"FE", x"FE", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"01", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"01", x"FF", x"01", x"FF", x"FC", x"02", x"00",
	x"00", x"FF", x"02", x"FD", x"01", x"FD", x"00", x"02", x"02", x"FF", x"00", x"FE",
	x"FE", x"01", x"01", x"00", x"FD", x"01", x"FF", x"FF", x"FE", x"FF", x"00", x"00",
	x"02", x"FC", x"FE", x"02", x"01", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FE",
	x"FF", x"01", x"FF", x"FD", x"FF", x"01", x"02", x"02", x"FC", x"FD", x"FE", x"02",
	x"00", x"FE", x"FE", x"01", x"02", x"02", x"FE", x"02", x"FF", x"FF", x"FF", x"FD",
	x"00", x"00", x"01", x"01", x"FE", x"02", x"FE", x"00", x"00", x"01", x"FF", x"00",
	x"FF", x"FE", x"FF", x"02", x"FF", x"FF", x"01", x"FE", x"01", x"02", x"FE", x"FF",
	x"FE", x"00", x"FE", x"00", x"FF", x"01", x"02", x"02", x"FE", x"01", x"FE", x"FD",
	x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"01", x"FE", x"01", x"FE", x"FE",
	x"00", x"02", x"00", x"01", x"02", x"00", x"00", x"FF", x"FD", x"FE", x"01", x"FF",
	x"01", x"01", x"01", x"FF", x"FE", x"FF", x"FE", x"00", x"00", x"FD", x"01", x"02",
	x"FE", x"FF", x"01", x"FE", x"00", x"00", x"00", x"FD", x"01", x"01", x"00", x"FE",
	x"FE", x"01", x"00", x"00", x"00", x"00", x"02", x"FF", x"00", x"FE", x"FE", x"00",
	x"FF", x"FD", x"02", x"00", x"03", x"FD", x"FE", x"FE", x"01", x"01", x"FE", x"FF",
	x"FF", x"04", x"00", x"FE", x"FD", x"FE", x"00", x"00", x"FF", x"FD", x"FE", x"05",
	x"01", x"FD", x"00", x"FF", x"01", x"FF", x"FE", x"FF", x"00", x"01", x"01", x"FE",
	x"FD", x"02", x"01", x"00", x"FE", x"00", x"FF", x"FF", x"FD", x"00", x"00", x"02",
	x"02", x"FC", x"FD", x"01", x"00", x"FF", x"01", x"FC", x"00", x"00", x"00", x"FD",
	x"FF", x"02", x"00", x"FE", x"00", x"FF", x"FF", x"00", x"FE", x"FF", x"FF", x"03",
	x"00", x"00", x"FE", x"FF", x"00", x"FD", x"FD", x"02", x"FF", x"01", x"02", x"FF",
	x"00", x"00", x"00", x"FD", x"FF", x"FE", x"01", x"01", x"02", x"FF", x"FF", x"00",
	x"FE", x"FE", x"FF", x"01", x"00", x"02", x"FF", x"FF", x"FE", x"FE", x"FE", x"02",
	x"00", x"00", x"03", x"FE", x"00", x"FF", x"FD", x"FF", x"00", x"00", x"FC", x"02",
	x"01", x"FF", x"FD", x"03", x"FF", x"FC", x"FF", x"01", x"FF", x"01", x"02", x"FF",
	x"FD", x"FD", x"00", x"FF", x"02", x"00", x"00", x"FD", x"00", x"00", x"FE", x"00",
	x"FE", x"00", x"01", x"03", x"FE", x"FE", x"00", x"FF", x"FD", x"FD", x"FF", x"00",
	x"02", x"02", x"FF", x"FC", x"FF", x"FF", x"00", x"FE", x"00", x"01", x"02", x"00",
	x"00", x"FF", x"FE", x"FF", x"FD", x"FF", x"03", x"01", x"00", x"00", x"FE", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"02", x"02", x"FF", x"FD", x"00", x"FF", x"00", x"FD",
	x"00", x"FE", x"03", x"FF", x"02", x"FE", x"01", x"01", x"FE", x"FE", x"FD", x"00",
	x"01", x"01", x"01", x"FF", x"01", x"00", x"FF", x"00", x"FF", x"00", x"01", x"FC",
	x"FE", x"00", x"03", x"FF", x"FF", x"FF", x"00", x"02", x"FF", x"FD", x"01", x"FF",
	x"00", x"00", x"FE", x"01", x"FE", x"01", x"FF", x"FD", x"00", x"00", x"FE", x"01",
	x"FE", x"01", x"FE", x"00", x"FF", x"FE", x"00", x"01", x"00", x"FF", x"01", x"00",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"00", x"FF", x"00", x"FE", x"FF",
	x"FF", x"FF", x"00", x"FF", x"01", x"00", x"FF", x"FE", x"00", x"01", x"00", x"FD",
	x"00", x"00", x"01", x"02", x"FF", x"01", x"FE", x"00", x"01", x"FE", x"FE", x"01",
	x"02", x"00", x"FE", x"00", x"FF", x"00", x"FE", x"FE", x"00", x"01", x"00", x"FE",
	x"02", x"FE", x"FE", x"01", x"FE", x"FE", x"03", x"00", x"00", x"FD", x"FE", x"00",
	x"01", x"01", x"FC", x"01", x"01", x"00", x"FF", x"FC", x"FF", x"FF", x"01", x"FF",
	x"00", x"03", x"00", x"FF", x"FE", x"FC", x"FE", x"01", x"FF", x"FF", x"02", x"01",
	x"01", x"00", x"FD", x"FE", x"FF", x"FE", x"FE", x"00", x"03", x"01", x"03", x"00",
	x"FC", x"FE", x"FF", x"FF", x"FF", x"00", x"FE", x"00", x"01", x"FF", x"00", x"00",
	x"00", x"FB", x"FF", x"00", x"00", x"01", x"02", x"FF", x"01", x"FD", x"FF", x"FD",
	x"00", x"01", x"FF", x"00", x"FE", x"01", x"01", x"03", x"FE", x"FF", x"FE", x"FD",
	x"00", x"01", x"04", x"00", x"00", x"00", x"FE", x"FF", x"FD", x"00", x"FE", x"00",
	x"01", x"00", x"00", x"00", x"01", x"FE", x"FE", x"FE", x"FE", x"FF", x"03", x"00",
	x"02", x"FF", x"FF", x"01", x"FE", x"00", x"00", x"00", x"FE", x"00", x"FE", x"00",
	x"00", x"00", x"FF", x"00", x"FE", x"FF", x"01", x"FF", x"01", x"FE", x"FE", x"FE",
	x"01", x"01", x"03", x"FF", x"FF", x"FC", x"FF", x"01", x"FF", x"FE", x"FE", x"00",
	x"01", x"00", x"FE", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"01", x"01", x"00",
	x"FE", x"FF", x"01", x"FF", x"00", x"01", x"00", x"00", x"FE", x"FE", x"FE", x"00",
	x"02", x"FF", x"01", x"FF", x"00", x"02", x"FE", x"00", x"FF", x"01", x"FF", x"FE",
	x"FD", x"00", x"00", x"02", x"FF", x"FF", x"FF", x"01", x"01", x"00", x"FF", x"FE",
	x"FF", x"00", x"00", x"FF", x"00", x"01", x"FD", x"FC", x"FD", x"00", x"01", x"00",
	x"FE", x"03", x"FE", x"00", x"FD", x"FF", x"FD", x"01", x"01", x"FF", x"FF", x"00",
	x"02", x"FE", x"FE", x"FC", x"FF", x"FF", x"01", x"00", x"01", x"01", x"FF", x"FF",
	x"FD", x"FE", x"01", x"00", x"00", x"01", x"00", x"01", x"FF", x"FE", x"FC", x"01",
	x"FF", x"FF", x"02", x"01", x"FF", x"00", x"FF", x"FD", x"FF", x"01", x"00", x"FE",
	x"03", x"FE", x"00", x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"FF", x"02", x"FF",
	x"FD", x"FE", x"FE", x"00", x"01", x"FF", x"FF", x"00", x"02", x"FE", x"FF", x"FC",
	x"00", x"FF", x"02", x"FE", x"00", x"00", x"00", x"FE", x"00", x"FE", x"00", x"01",
	x"FF", x"00", x"00", x"00", x"01", x"FE", x"FF", x"FF", x"FF", x"00", x"02", x"00",
	x"00", x"00", x"FE", x"FE", x"00", x"02", x"00", x"FD", x"00", x"FE", x"01", x"01",
	x"FE", x"FF", x"FF", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FE", x"01",
	x"01", x"01", x"FE", x"FE", x"FF", x"00", x"FD", x"FF", x"00", x"FF", x"02", x"01",
	x"00", x"FE", x"00", x"00", x"FC", x"FF", x"FF", x"02", x"01", x"00", x"00", x"FF",
	x"FF", x"FF", x"FE", x"00", x"00", x"00", x"00", x"FF", x"FE", x"02", x"FE", x"00",
	x"FE", x"FF", x"00", x"01", x"FE", x"FE", x"00", x"FF", x"01", x"FC", x"01", x"FF",
	x"02", x"01", x"FD", x"FE", x"FF", x"00", x"00", x"FF", x"FE", x"02", x"FE", x"01",
	x"00", x"01", x"FE", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FE", x"02", x"FF",
	x"FF", x"00", x"FF", x"FF", x"02", x"FE", x"FE", x"FE", x"02", x"01", x"FD", x"00",
	x"FF", x"01", x"02", x"00", x"FC", x"00", x"FE", x"00", x"FD", x"FF", x"00", x"03",
	x"01", x"01", x"FD", x"FE", x"FD", x"02", x"FF", x"01", x"03", x"FE", x"00", x"FE",
	x"00", x"FF", x"FF", x"FE", x"FD", x"02", x"01", x"00", x"00", x"03", x"FE", x"FE",
	x"FD", x"01", x"FE", x"03", x"FF", x"FF", x"FE", x"01", x"01", x"FF", x"FE", x"FF",
	x"FE", x"01", x"00", x"00", x"FF", x"01", x"00", x"FF", x"FF", x"FE", x"00", x"01",
	x"FF", x"00", x"FE", x"01", x"FF", x"02", x"FF", x"01", x"FC", x"FF", x"01", x"00",
	x"00", x"FF", x"01", x"FF", x"00", x"FF", x"FF", x"FE", x"01", x"01", x"FF", x"FF",
	x"FF", x"FF", x"02", x"00", x"FE", x"FE", x"FF", x"01", x"00", x"00", x"00", x"FF",
	x"FF", x"FE", x"FE", x"00", x"00", x"FD", x"01", x"02", x"00", x"FE", x"00", x"FF",
	x"00", x"FF", x"FF", x"FE", x"00", x"00", x"00", x"FE", x"00", x"FE", x"01", x"FF",
	x"FF", x"FF", x"00", x"01", x"FF", x"00", x"FF", x"FD", x"FF", x"03", x"FF", x"00",
	x"FE", x"FE", x"00", x"FF", x"01", x"FC", x"01", x"00", x"01", x"FE", x"00", x"FF",
	x"FE", x"00", x"00", x"FF", x"00", x"01", x"01", x"00", x"FF", x"FE", x"00", x"FE",
	x"01", x"FF", x"00", x"01", x"00", x"01", x"FF", x"00", x"00", x"FD", x"FE", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"FE", x"00", x"FD", x"02", x"FF", x"01", x"01",
	x"FD", x"00", x"FE", x"01", x"FE", x"FF", x"FF", x"FF", x"FF", x"01", x"00", x"02",
	x"01", x"FE", x"FE", x"FD", x"FF", x"01", x"01", x"01", x"FF", x"02", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"00", x"FE", x"00", x"01", x"00", x"01", x"FE", x"FE",
	x"FF", x"00", x"FF", x"01", x"00", x"FD", x"00", x"02", x"00", x"FE", x"00", x"FE",
	x"FE", x"00", x"01", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"01", x"00", x"FE", x"FE", x"00", x"FF", x"00", x"FF", x"FE", x"00", x"00",
	x"03", x"FE", x"FE", x"FD", x"01", x"01", x"00", x"FD", x"FE", x"00", x"00", x"00",
	x"FE", x"00", x"00", x"01", x"FF", x"FD", x"FE", x"00", x"03", x"01", x"FF", x"01",
	x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"01", x"FF", x"00", x"FF", x"FD",
	x"00", x"FE", x"02", x"FF", x"02", x"00", x"00", x"02", x"FC", x"FD", x"FD", x"01",
	x"01", x"FF", x"00", x"01", x"00", x"02", x"FF", x"FD", x"FE", x"01", x"FF", x"FE",
	x"00", x"01", x"02", x"01", x"FE", x"FE", x"FD", x"FF", x"01", x"FF", x"FE", x"00",
	x"00", x"00", x"FE", x"01", x"00", x"00", x"00", x"01", x"FC", x"00", x"FE", x"00",
	x"FE", x"01", x"FE", x"00", x"00", x"FE", x"02", x"00", x"00", x"FD", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"FF", x"01", x"FE", x"01", x"FD", x"01", x"FF", x"FE",
	x"FE", x"00", x"00", x"FF", x"00", x"01", x"FF", x"FF", x"01", x"FE", x"FF", x"FC",
	x"00", x"FE", x"02", x"01", x"00", x"FD", x"01", x"01", x"00", x"FE", x"FD", x"FF",
	x"02", x"FF", x"01", x"FE", x"FF", x"00", x"01", x"FE", x"FE", x"02", x"02", x"00",
	x"FE", x"FF", x"00", x"01", x"FF", x"FD", x"FF", x"00", x"02", x"FE", x"00", x"FF",
	x"00", x"FF", x"FD", x"00", x"00", x"02", x"00", x"FF", x"02", x"01", x"FF", x"00",
	x"FE", x"FE", x"01", x"01", x"00", x"FE", x"00", x"02", x"00", x"FF", x"FE", x"FF",
	x"00", x"01", x"FD", x"FF", x"00", x"03", x"FF", x"FD", x"FE", x"01", x"00", x"FF",
	x"00", x"FE", x"00", x"00", x"FE", x"FE", x"01", x"01", x"02", x"FD", x"FF", x"FF",
	x"00", x"01", x"FF", x"FD", x"FF", x"00", x"01", x"00", x"FF", x"FF", x"01", x"FE",
	x"FF", x"00", x"FF", x"FF", x"00", x"01", x"FE", x"01", x"00", x"FE", x"01", x"FD",
	x"01", x"FF", x"01", x"FE", x"01", x"02", x"FF", x"FE", x"FF", x"FF", x"00", x"01",
	x"00", x"FF", x"FF", x"01", x"FF", x"FF", x"FD", x"FE", x"01", x"FF", x"00", x"01",
	x"FF", x"01", x"FF", x"00", x"FD", x"FE", x"00", x"02", x"FD", x"00", x"FF", x"FE",
	x"01", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"01", x"FF", x"02", x"FE", x"02",
	x"FE", x"FF", x"00", x"FF", x"FE", x"01", x"FF", x"FF", x"00", x"FF", x"00", x"02",
	x"FF", x"00", x"FE", x"FF", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"01",
	x"FF", x"00", x"00", x"00", x"FE", x"00", x"00", x"00", x"FF", x"00", x"FC", x"FF",
	x"02", x"01", x"FE", x"00", x"00", x"FF", x"FF", x"FF", x"FD", x"00", x"00", x"FF",
	x"FF", x"01", x"02", x"01", x"FF", x"FC", x"FE", x"00", x"00", x"FF", x"01", x"FF",
	x"00", x"02", x"FD", x"FF", x"FF", x"00", x"FF", x"FD", x"00", x"00", x"01", x"01",
	x"01", x"FD", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FE", x"FE", x"FF",
	x"02", x"FF", x"00", x"FD", x"00", x"01", x"00", x"00", x"FE", x"00", x"01", x"FF",
	x"FD", x"FE", x"00", x"03", x"FE", x"00", x"FF", x"00", x"00", x"FE", x"01", x"FD",
	x"00", x"FE", x"01", x"FF", x"01", x"00", x"FF", x"FE", x"00", x"FD", x"00", x"00",
	x"00", x"FE", x"01", x"00", x"00", x"FE", x"00", x"01", x"00", x"FF", x"FE", x"FE",
	x"01", x"01", x"01", x"FD", x"FF", x"FF", x"FF", x"FF", x"00", x"FE", x"01", x"FF",
	x"01", x"FE", x"FF", x"00", x"FF", x"02", x"00", x"FF", x"FF", x"02", x"FF", x"FF",
	x"FE", x"FF", x"00", x"01", x"00", x"FF", x"00", x"FE", x"03", x"FD", x"00", x"FF",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"02", x"FF", x"FF", x"01", x"FE", x"FE",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"02", x"FF", x"00", x"FE", x"01",
	x"00", x"FF", x"FF", x"FE", x"03", x"FF", x"01", x"FD", x"FF", x"FD", x"03", x"FE",
	x"FE", x"FE", x"01", x"01", x"FF", x"00", x"FE", x"03", x"00", x"00", x"FD", x"FE",
	x"00", x"FF", x"00", x"FD", x"01", x"FF", x"01", x"FE", x"FF", x"00", x"02", x"FE",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"01", x"FF", x"FF", x"FF", x"01",
	x"FF", x"00", x"FD", x"FF", x"00", x"02", x"FF", x"FE", x"FE", x"02", x"01", x"FF",
	x"FE", x"FF", x"00", x"00", x"01", x"FE", x"FE", x"00", x"01", x"FF", x"FE", x"01",
	x"FF", x"FF", x"00", x"FE", x"FF", x"FF", x"FF", x"01", x"FE", x"02", x"FE", x"00",
	x"00", x"01", x"FF", x"FD", x"FD", x"00", x"FF", x"01", x"00", x"01", x"FE", x"02",
	x"00", x"FF", x"FD", x"00", x"FE", x"01", x"00", x"00", x"01", x"00", x"FF", x"FF",
	x"FF", x"01", x"00", x"00", x"FF", x"00", x"FF", x"02", x"FE", x"FF", x"FF", x"00",
	x"FF", x"FF", x"00", x"02", x"FF", x"FE", x"FF", x"00", x"FE", x"01", x"FF", x"01",
	x"FE", x"00", x"FE", x"01", x"FF", x"00", x"01", x"FF", x"FF", x"FE", x"00", x"00",
	x"00", x"FF", x"02", x"01", x"FE", x"FD", x"01", x"FF", x"00", x"FF", x"01", x"FF",
	x"02", x"00", x"00", x"FB", x"01", x"00", x"FF", x"FF", x"00", x"01", x"FF", x"01",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"01", x"FE", x"FF", x"FE",
	x"00", x"FD", x"FF", x"FF", x"03", x"01", x"FF", x"FE", x"00", x"FE", x"01", x"FE",
	x"FE", x"FF", x"02", x"01", x"FE", x"00", x"FE", x"00", x"00", x"00", x"FE", x"01",
	x"01", x"00", x"00", x"FE", x"FE", x"FF", x"FF", x"FF", x"01", x"01", x"FE", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FE", x"01", x"00", x"00", x"FF", x"FF", x"00",
	x"FF", x"01", x"FD", x"01", x"FE", x"01", x"00", x"FE", x"FE", x"00", x"01", x"FF",
	x"00", x"FF", x"01", x"FF", x"03", x"FD", x"00", x"FE", x"00", x"FF", x"00", x"FF",
	x"00", x"FE", x"00", x"FE", x"00", x"00", x"FF", x"00", x"01", x"00", x"00", x"00",
	x"FD", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FE", x"00", x"FF", x"00", x"FD",
	x"02", x"FF", x"00", x"00", x"FF", x"02", x"FF", x"FF", x"FF", x"00", x"FD", x"FF",
	x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"01", x"01", x"FE", x"01", x"FE",
	x"FD", x"01", x"FF", x"00", x"00", x"00", x"00", x"00", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"FF", x"02", x"FF", x"FF", x"FE", x"FF", x"FD", x"00",
	x"01", x"01", x"00", x"00", x"FE", x"00", x"FF", x"FF", x"00", x"00", x"FE", x"01",
	x"FE", x"00", x"FF", x"FF", x"00", x"00", x"FE", x"01", x"00", x"02", x"FE", x"01",
	x"FD", x"FF", x"FE", x"02", x"FF", x"FF", x"00", x"00", x"FF", x"02", x"00", x"FE",
	x"00", x"00", x"FE", x"00", x"FE", x"02", x"FF", x"01", x"FF", x"FF", x"01", x"00",
	x"00", x"FF", x"FE", x"FE", x"00", x"00", x"FF", x"02", x"00", x"FF", x"FE", x"FF",
	x"00", x"00", x"01", x"00", x"01", x"00", x"FF", x"FE", x"FF", x"FE", x"01", x"FF",
	x"01", x"00", x"00", x"01", x"FF", x"FE", x"FE", x"FF", x"FF", x"01", x"FE", x"01",
	x"01", x"00", x"FF", x"FE", x"00", x"FE", x"01", x"FE", x"FE", x"01", x"01", x"00",
	x"FF", x"01", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"01", x"00", x"00", x"FE",
	x"00", x"00", x"FF", x"FE", x"FF", x"01", x"00", x"00", x"FF", x"02", x"FE", x"FE",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"FF", x"01", x"FD", x"FF", x"FE",
	x"FF", x"FF", x"00", x"02", x"FF", x"01", x"00", x"FE", x"FD", x"FF", x"FF", x"01",
	x"01", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FD", x"01", x"FF", x"01", x"00",
	x"FF", x"01", x"00", x"01", x"FF", x"FC", x"01", x"FF", x"01", x"00", x"FE", x"FF",
	x"00", x"00", x"FF", x"FF", x"01", x"01", x"FE", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FE", x"01", x"00", x"FF", x"FC", x"01", x"00", x"00", x"FE", x"00", x"02",
	x"FF", x"00", x"FD", x"FD", x"01", x"00", x"00", x"FE", x"01", x"01", x"FF", x"FE",
	x"FF", x"FF", x"01", x"FF", x"FF", x"FD", x"00", x"00", x"FF", x"FE", x"00", x"00",
	x"01", x"FF", x"00", x"FE", x"00", x"FF", x"FF", x"FE", x"00", x"00", x"01", x"00",
	x"FF", x"FF", x"FE", x"00", x"FF", x"01", x"FE", x"02", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"00", x"00", x"00", x"01", x"FF", x"00", x"00", x"00", x"00", x"FD", x"FF",
	x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"01",
	x"00", x"00", x"00", x"FF", x"FE", x"00", x"FE", x"FF", x"00", x"00", x"00", x"00",
	x"01", x"FF", x"FD", x"FF", x"01", x"00", x"FF", x"FF", x"FF", x"01", x"00", x"FF",
	x"FD", x"00", x"FF", x"02", x"FE", x"00", x"FF", x"01", x"00", x"00", x"FF", x"00",
	x"00", x"FF", x"FE", x"FE", x"02", x"00", x"FF", x"FE", x"FF", x"00", x"00", x"00",
	x"FE", x"00", x"00", x"00", x"FF", x"FF", x"01", x"FF", x"00", x"FF", x"FE", x"FE",
	x"02", x"01", x"FE", x"FE", x"01", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FE",
	x"FF", x"FF", x"01", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"00", x"00",
	x"FF", x"01", x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"FF",
	x"01", x"FE", x"00", x"00", x"FE", x"FE", x"FE", x"01", x"01", x"00", x"FF", x"00",
	x"00", x"FF", x"00", x"00", x"FE", x"00", x"00", x"FF", x"01", x"FF", x"01", x"FF",
	x"00", x"FE", x"FE", x"00", x"01", x"FF", x"FF", x"FF", x"02", x"FF", x"01", x"FE",
	x"00", x"FE", x"01", x"FF", x"FF", x"01", x"01", x"FF", x"FF", x"FF", x"FE", x"00",
	x"01", x"FE", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"00",
	x"00", x"03", x"00", x"FF", x"FE", x"00", x"FF", x"FF", x"00", x"FE", x"02", x"00",
	x"01", x"FF", x"FD", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"02", x"02", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"FE", x"00", x"00",
	x"FE", x"00", x"FF", x"FF", x"02", x"00", x"00", x"00", x"FF", x"FE", x"00", x"FF",
	x"01", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"01", x"01", x"00", x"FE", x"00",
	x"01", x"00", x"FF", x"FE", x"FD", x"02", x"00", x"FF", x"00", x"FE", x"00", x"FF",
	x"00", x"FD", x"01", x"01", x"01", x"00", x"FE", x"01", x"FE", x"00", x"FE", x"FE",
	x"00", x"02", x"FF", x"FF", x"FE", x"01", x"FF", x"FF", x"00", x"01", x"02", x"FF",
	x"FE", x"FE", x"FF", x"01", x"00", x"FE", x"FE", x"00", x"01", x"00", x"FF", x"FE",
	x"00", x"00", x"00", x"FF", x"FD", x"02", x"FF", x"00", x"FE", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"FE", x"00", x"FF", x"00", x"00", x"00", x"FF",
	x"00", x"FE", x"00", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"01", x"FF",
	x"00", x"FD", x"00", x"FF", x"01", x"FF", x"00", x"FF", x"FF", x"FE", x"01", x"FE",
	x"00", x"00", x"00", x"00", x"FD", x"00", x"FF", x"01", x"FF", x"FE", x"FE", x"00",
	x"02", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"00", x"FF", x"FF", x"01", x"FF",
	x"FC", x"00", x"01", x"01", x"00", x"FF", x"FE", x"FF", x"00", x"01", x"FC", x"01",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"00", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"01", x"FF", x"FE", x"FF", x"01", x"00", x"00", x"FF", x"FE", x"FF",
	x"02", x"00", x"FE", x"00", x"00", x"01", x"FE", x"FE", x"FE", x"00", x"01", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"01", x"01", x"00", x"FF",
	x"00", x"FF", x"FE", x"00", x"FF", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"01", x"03", x"FE", x"00", x"FD", x"FF", x"FE",
	x"01", x"00", x"00", x"01", x"00", x"FE", x"FE", x"00", x"FE", x"00", x"FF", x"00",
	x"00", x"00", x"01", x"FF", x"FF", x"FF", x"00", x"FE", x"01", x"FE", x"02", x"FF",
	x"FE", x"00", x"00", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"FE", x"FF", x"00",
	x"00", x"01", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"03", x"FF", x"00",
	x"FE", x"FD", x"FF", x"00", x"01", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"FE", x"FF", x"00", x"00", x"FF", x"02", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"FF", x"01",
	x"01", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FD", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"FF", x"00",
	x"00", x"00", x"FF", x"FE", x"00", x"FF", x"FF", x"01", x"FE", x"00", x"00", x"00",
	x"00", x"00", x"01", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"01", x"00",
	x"FE", x"00", x"FF", x"00", x"FE", x"01", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"01", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"01", x"FF", x"00", x"01", x"FF", x"FF", x"FF", x"00",
	x"FE", x"00", x"FE", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE",
	x"FF", x"FF", x"FF", x"01", x"FE", x"01", x"FD", x"00", x"FE", x"01", x"FE", x"FF",
	x"FF", x"FF", x"00", x"FE", x"FF", x"00", x"FE", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"FE", x"FF", x"01", x"00", x"FF", x"00", x"01", x"FF",
	x"01", x"00", x"FE", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"01", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"FE", x"FF", x"01", x"00", x"00", x"FE", x"FE",
	x"00", x"00", x"00", x"FD", x"01", x"00", x"00", x"FE", x"01", x"FF", x"FE", x"FF",
	x"00", x"00", x"00", x"01", x"FE", x"FE", x"00", x"00", x"FF", x"FF", x"00", x"01",
	x"00", x"01", x"FE", x"FE", x"00", x"00", x"00", x"00", x"FF", x"00", x"01", x"FF",
	x"FE", x"FF", x"00", x"00", x"FE", x"FF", x"00", x"02", x"00", x"00", x"FE", x"00",
	x"FE", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00",
	x"FF", x"FE", x"00", x"00", x"00", x"02", x"FF", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"FE", x"00", x"00", x"00", x"01", x"FE", x"FF", x"FF", x"00", x"FE", x"00",
	x"00", x"FF", x"02", x"FE", x"FF", x"FD", x"00", x"FF", x"00", x"00", x"00", x"FE",
	x"FF", x"01", x"00", x"00", x"FD", x"FF", x"00", x"00", x"00", x"FF", x"01", x"00",
	x"01", x"FC", x"FE", x"FF", x"00", x"FF", x"01", x"FE", x"00", x"00", x"01", x"FF",
	x"FF", x"00", x"00", x"FD", x"00", x"01", x"FF", x"01", x"FF", x"FF", x"FF", x"00",
	x"02", x"FD", x"FF", x"FF", x"00", x"FE", x"FD", x"01", x"00", x"01", x"00", x"FE",
	x"FE", x"00", x"00", x"FE", x"00", x"00", x"00", x"FF", x"00", x"FE", x"01", x"FF",
	x"FF", x"FF", x"FE", x"00", x"FE", x"02", x"FE", x"FF", x"FF", x"01", x"FF", x"FF",
	x"00", x"01", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"01", x"FF", x"01",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FE", x"00", x"FF", x"FF", x"FF", x"01", x"FF", x"00", x"FF", x"00", x"01",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"01", x"FE",
	x"00", x"FE", x"FF", x"00", x"01", x"FF", x"FE", x"FF", x"01", x"FF", x"FF", x"FF",
	x"01", x"FF", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"01",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FE", x"00", x"FE",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"FE", x"00", x"00", x"FF",
	x"00", x"FF", x"01", x"00", x"01", x"FF", x"FF", x"FE", x"01", x"FF", x"00", x"FF",
	x"FF", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00",
	x"FF", x"FE", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FE", x"01", x"FE", x"01",
	x"FE", x"01", x"FE", x"FF", x"00", x"FF", x"FF", x"01", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FE", x"01", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"00", x"01", x"FF", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FD", x"01", x"01",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FE", x"01", x"FD", x"01", x"FE", x"01", x"01", x"FE", x"00",
	x"FF", x"00", x"01", x"FF", x"00", x"FE", x"00", x"00", x"00", x"FE", x"00", x"FD",
	x"01", x"00", x"00", x"FF", x"FE", x"03", x"FF", x"00", x"FE", x"FF", x"01", x"FE",
	x"FF", x"FE", x"01", x"FF", x"01", x"00", x"FF", x"FE", x"00", x"00", x"01", x"FF",
	x"FE", x"00", x"FF", x"01", x"00", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"01",
	x"FE", x"FF", x"FE", x"01", x"FE", x"00", x"FF", x"01", x"FF", x"FE", x"00", x"00",
	x"FF", x"01", x"FE", x"01", x"FE", x"00", x"00", x"00", x"FF", x"01", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"FE", x"00", x"FE", x"FF", x"00", x"02", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"01", x"01", x"01", x"FF", x"00",
	x"00", x"01", x"FD", x"FF", x"FE", x"00", x"00", x"00", x"00", x"FE", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FE", x"01", x"FF", x"FE", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"01", x"FF", x"00", x"FE", x"00", x"00", x"FF", x"00",
	x"FE", x"FF", x"01", x"00", x"02", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF",
	x"01", x"00", x"00", x"FE", x"FF", x"FF", x"FF", x"01", x"FE", x"FE", x"00", x"01",
	x"03", x"FE", x"00", x"FD", x"FF", x"01", x"FE", x"00", x"FE", x"01", x"00", x"00",
	x"FD", x"00", x"FE", x"01", x"FF", x"FF", x"01", x"FF", x"00", x"FF", x"FE", x"00",
	x"FF", x"00", x"01", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"01", x"00", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE",
	x"01", x"FD", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"FE", x"FF",
	x"FE", x"FF", x"00", x"FE", x"01", x"FF", x"01", x"FF", x"01", x"FF", x"00", x"FF",
	x"FF", x"FF", x"01", x"FF", x"00", x"00", x"01", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"01", x"00", x"FE", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"FE", x"00", x"00", x"FE", x"00", x"00", x"00", x"FE", x"00", x"FF", x"01",
	x"FF", x"FF", x"01", x"FE", x"01", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FE",
	x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"01", x"FD", x"00", x"FE", x"00",
	x"00", x"FE", x"00", x"00", x"FF", x"00", x"FE", x"01", x"00", x"FF", x"FF", x"FE",
	x"00", x"FF", x"01", x"FF", x"00", x"00", x"00", x"FF", x"01", x"FF", x"00", x"FF",
	x"FF", x"00", x"FD", x"00", x"01", x"01", x"01", x"FF", x"01", x"FF", x"00", x"FF",
	x"FF", x"01", x"FF", x"FF", x"01", x"FD", x"02", x"FF", x"01", x"00", x"FE", x"FE",
	x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"00", x"01", x"FF", x"00", x"FF", x"00", x"FE", x"00", x"FE", x"01", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"01", x"01", x"00",
	x"FE", x"00", x"FE", x"00", x"FF", x"FE", x"00", x"01", x"01", x"FF", x"FE", x"FF",
	x"00", x"00", x"00", x"FE", x"FF", x"00", x"01", x"FF", x"00", x"00", x"FF", x"01",
	x"FD", x"FF", x"FF", x"01", x"FF", x"FF", x"FE", x"FF", x"FF", x"01", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FE", x"00", x"00", x"02", x"00",
	x"FF", x"FF", x"00", x"00", x"FF", x"FE", x"FF", x"00", x"01", x"00", x"FE", x"FF",
	x"01", x"01", x"FF", x"FD", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"00", x"02", x"FE", x"FF", x"FF", x"01", x"FE", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FF", x"00", x"01", x"FF",
	x"01", x"FE", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"01", x"FF", x"00",
	x"00", x"00", x"FE", x"01", x"FF", x"01", x"00", x"FE", x"01", x"FE", x"00", x"FE",
	x"FF", x"FF", x"FF", x"01", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FE", x"02", x"FF", x"01", x"FE", x"FE", x"FF", x"00", x"FF", x"01", x"FF", x"FF",
	x"00", x"00", x"01", x"00", x"00", x"01", x"FF", x"FF", x"FE", x"FE", x"01", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"01", x"00", x"FF", x"FF", x"FF", x"01", x"FF", x"FF", x"01", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"02", x"FE", x"00", x"FE", x"01", x"00", x"01", x"FF", x"FE",
	x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"00", x"00",
	x"FF", x"00", x"00", x"FF", x"01", x"FE", x"FF", x"01", x"00", x"01", x"00", x"FF",
	x"00", x"FF", x"00", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF",
	x"01", x"FE", x"00", x"00", x"FF", x"01", x"FE", x"00", x"00", x"00", x"FE", x"00",
	x"FF", x"00", x"FF", x"02", x"FE", x"FE", x"00", x"00", x"FE", x"01", x"00", x"01",
	x"00", x"FF", x"FE", x"00", x"00", x"00", x"FF", x"00", x"02", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FE", x"00", x"FF", x"00", x"FF", x"01", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"FE", x"00", x"FF", x"00",
	x"00", x"FF", x"00", x"FF", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"00", x"FF", x"01", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FE", x"00", x"FE", x"01", x"FE", x"02", x"01", x"FF", x"00",
	x"FD", x"00", x"00", x"FD", x"01", x"00", x"00", x"01", x"FF", x"FF", x"FF", x"FF",
	x"01", x"00", x"00", x"FE", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"01", x"FE", x"01", x"FF", x"FF", x"FF", x"01", x"FE", x"00", x"01", x"FF", x"FF",
	x"FF", x"01", x"FE", x"01", x"FD", x"00", x"FE", x"00", x"00", x"00", x"01", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"01", x"FF", x"FD", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"01",
	x"FE", x"00", x"FF", x"00", x"FF", x"01", x"FF", x"FF", x"01", x"01", x"FE", x"FF",
	x"FF", x"00", x"02", x"FE", x"00", x"FF", x"00", x"FF", x"FD", x"01", x"FF", x"01",
	x"00", x"00", x"FE", x"00", x"FE", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"FE",
	x"01", x"00", x"00", x"FE", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"FE", x"FF", x"FF", x"02", x"00", x"00", x"FE", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"01", x"01", x"00", x"00", x"FD", x"01", x"00", x"01", x"FF", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"00", x"FE", x"01", x"FE", x"01", x"FF", x"01", x"00",
	x"FE", x"FE", x"01", x"00", x"00", x"00", x"FF", x"FF", x"01", x"FE", x"FF", x"FD",
	x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"01", x"FF", x"00", x"FF", x"00", x"FD", x"00", x"00",
	x"00", x"00", x"FE", x"FE", x"00", x"01", x"01", x"FE", x"00", x"FE", x"01", x"FF",
	x"FF", x"FE", x"01", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FE",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FF",
	x"01", x"00", x"FF", x"00", x"FE", x"00", x"00", x"00", x"FE", x"00", x"FF", x"00",
	x"00", x"FF", x"FE", x"FF", x"01", x"FF", x"00", x"01", x"FF", x"00", x"00", x"01",
	x"FE", x"FF", x"00", x"FF", x"00", x"00", x"FE", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00",
	x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"00", x"FF", x"01", x"FF", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"01", x"FE", x"00", x"FF",
	x"01", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"01", x"FF",
	x"FF", x"FF", x"FE", x"00", x"FE", x"00", x"FE", x"01", x"FF", x"00", x"FF", x"00",
	x"FF", x"01", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"01", x"00", x"FF", x"FE", x"00", x"FE", x"01", x"FF", x"FF", x"00", x"FF",
	x"00", x"FE", x"00", x"FE", x"00", x"00", x"00", x"00", x"FF", x"00", x"01", x"FF",
	x"FE", x"FE", x"FF", x"02", x"00", x"00", x"FF", x"FF", x"00", x"FE", x"00", x"FF",
	x"FF", x"01", x"FF", x"00", x"FF", x"00", x"01", x"FF", x"00", x"FF", x"FF", x"FF",
	x"01", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FE", x"FE",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"FE", x"00", x"FE", x"00", x"FF", x"00",
	x"00", x"FF", x"00", x"FF", x"02", x"FF", x"FF", x"FE", x"00", x"01", x"FF", x"FF",
	x"00", x"00", x"01", x"FF", x"FE", x"FE", x"01", x"00", x"FF", x"FE", x"FF", x"00",
	x"FF", x"01", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"01", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"FD", x"00", x"01", x"FF", x"00", x"FE", x"00",
	x"FF", x"FF", x"01", x"FE", x"01", x"FE", x"01", x"00", x"FF", x"FE", x"FF", x"FF",
	x"00", x"FF", x"01", x"00", x"00", x"00", x"FE", x"01", x"FE", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"01", x"00", x"00", x"00",
	x"00", x"FF", x"01", x"00", x"00", x"FF", x"02", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"FF", x"00", x"FF", x"01", x"FF", x"FF", x"FF", x"00", x"01", x"FE", x"00",
	x"FF", x"FF", x"FE", x"00", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"01", x"00",
	x"FF", x"FF", x"FE", x"01", x"01", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FE",
	x"00", x"FF", x"01", x"00", x"FF", x"00", x"FF", x"FE", x"01", x"FE", x"00", x"00",
	x"01", x"01", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"01", x"01", x"01",
	x"FF", x"00", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"FF", x"01", x"00", x"FF",
	x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"FF", x"FF", x"FE", x"00",
	x"00", x"01", x"FF", x"FE", x"00", x"FF", x"01", x"FF", x"01", x"FF", x"FF", x"FF",
	x"00", x"FD", x"00", x"00", x"00", x"00", x"FE", x"00", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"00",
	x"00", x"FF", x"00", x"01", x"FE", x"FE", x"01", x"00", x"00", x"FE", x"FE", x"FF",
	x"00", x"00", x"01", x"FE", x"01", x"FE", x"00", x"FE", x"FF", x"FF", x"01", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"FE", x"00", x"FF", x"00", x"FE", x"01", x"FF",
	x"00", x"00", x"FF", x"00", x"FE", x"00", x"FF", x"01", x"00", x"00", x"FE", x"00",
	x"FE", x"01", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FE", x"00",
	x"FF", x"FF", x"00", x"00", x"01", x"FE", x"01", x"FE", x"00", x"FF", x"FF", x"FF",
	x"01", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"01", x"FD", x"00", x"FF", x"01",
	x"FF", x"FF", x"01", x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"00", x"00", x"FF", x"01", x"00", x"FF",
	x"FF", x"00", x"FE", x"00", x"FF", x"01", x"00", x"FE", x"00", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"02", x"FF", x"01", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FE", x"01", x"00", x"00",
	x"FE", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FE", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"01", x"00",
	x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF",
	x"FE", x"00", x"00", x"FF", x"00", x"FF", x"00", x"01", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FE", x"00", x"00", x"01", x"FE", x"FF", x"00", x"00", x"00", x"FD",
	x"00", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"02", x"FE", x"01", x"FE", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FE", x"00", x"00", x"FE", x"FF", x"FE", x"01", x"01",
	x"00", x"01", x"FF", x"FF", x"01", x"FE", x"FF", x"00", x"FF", x"01", x"FF", x"01",
	x"FF", x"00", x"FF", x"FF", x"FE", x"01", x"FF", x"00", x"FF", x"01", x"FE", x"00",
	x"FF", x"FF", x"02", x"FE", x"FF", x"00", x"FF", x"01", x"FF", x"00", x"FF", x"FF",
	x"01", x"FE", x"00", x"FE", x"FF", x"01", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"01", x"FE",
	x"00", x"FF", x"00", x"FE", x"00", x"FF", x"00", x"FF", x"01", x"FF", x"00", x"FE",
	x"FF", x"FF", x"01", x"FF", x"00", x"00", x"00", x"FE", x"00", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"01", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"01", x"FF", x"01", x"FE", x"FE", x"01", x"FF", x"01", x"FF", x"00", x"00", x"FE",
	x"FF", x"FF", x"FF", x"01", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"FF",
	x"FF", x"00", x"FF", x"00", x"01", x"FF", x"00", x"FE", x"00", x"FD", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"FF", x"00", x"00", x"FE", x"FF",
	x"00", x"00", x"01", x"FE", x"01", x"FE", x"FF", x"01", x"00", x"FF", x"FF", x"01",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"01", x"FE", x"00",
	x"FF", x"FF", x"00", x"02", x"FF", x"FF", x"FF", x"FE", x"01", x"FF", x"00", x"00",
	x"00", x"00", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"01",
	x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FE", x"FF", x"FF", x"01", x"00", x"00",
	x"FF", x"FF", x"01", x"FF", x"FE", x"FF", x"00", x"FF", x"01", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"01", x"FF", x"FF", x"FF", x"01", x"FE",
	x"FF", x"00", x"FF", x"FF", x"FE", x"00", x"FF", x"01", x"FE", x"00", x"FF", x"01",
	x"FE", x"FF", x"FE", x"01", x"FF", x"FF", x"00", x"00", x"00", x"FE", x"01", x"FE",
	x"00", x"00", x"00", x"FF", x"01", x"FF", x"FF", x"FF", x"01", x"FF", x"FF", x"FF",
	x"00", x"01", x"FF", x"00", x"FD", x"FF", x"00", x"00", x"00", x"FE", x"FF", x"01",
	x"00", x"FF", x"FF", x"FF", x"00", x"FE", x"00", x"00", x"00", x"01", x"00", x"FE",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FE", x"00", x"FF",
	x"00", x"FE", x"01", x"FE", x"00", x"FF", x"FE", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"01", x"FF", x"FF", x"FF", x"FE", x"01", x"00", x"00", x"FE", x"00", x"01",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"02", x"FF", x"FF",
	x"FF", x"FF", x"00", x"01", x"00", x"FF", x"FE", x"01", x"FE", x"01", x"FF", x"FF",
	x"00", x"01", x"00", x"FF", x"FE", x"00", x"FF", x"01", x"FE", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FE", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"01",
	x"FF", x"FD", x"00", x"00", x"02", x"FF", x"FF", x"00", x"01", x"FF", x"FF", x"FE",
	x"01", x"01", x"FF", x"FF", x"FE", x"01", x"00", x"00", x"FE", x"FE", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"01", x"FF", x"FE", x"00", x"00", x"00", x"00", x"00",
	x"00", x"01", x"FE", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"02", x"FF",
	x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"01", x"FF", x"00", x"FE",
	x"FF", x"00", x"00", x"FF", x"FF", x"01", x"FF", x"00", x"FE", x"00", x"00", x"00",
	x"00", x"FE", x"00", x"00", x"00", x"00", x"FF", x"00", x"FE", x"00", x"00", x"FF",
	x"FF", x"FE", x"FF", x"00", x"00", x"FE", x"00", x"FF", x"01", x"00", x"00", x"FE",
	x"01", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"01", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"01", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"01", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"01", x"FF", x"01", x"FD", x"FF", x"FF", x"01", x"00", x"FF", x"FF", x"FF", x"01",
	x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"01", x"FE", x"00", x"00", x"00", x"FE",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"00", x"FF",
	x"01", x"00", x"00", x"FE", x"01", x"FF", x"FE", x"FF", x"FF", x"01", x"FF", x"00",
	x"FF", x"FE", x"00", x"00", x"00", x"FE", x"01", x"FF", x"00", x"FE", x"01", x"00",
	x"00", x"00", x"FE", x"00", x"00", x"01", x"FF", x"FE", x"01", x"00", x"01", x"FF",
	x"00", x"FF", x"01", x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"01", x"FF", x"FE", x"01", x"FF", x"FF", x"00",
	x"FD", x"01", x"00", x"01", x"FE", x"00", x"00", x"FF", x"FE", x"00", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"02", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"01", x"00",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"01",
	x"00", x"FF", x"FE", x"FF", x"01", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"01", x"FF", x"FF", x"00", x"FF", x"01", x"00", x"FE", x"00",
	x"FF", x"00", x"FE", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"01", x"FF", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FF", x"01", x"FF", x"00", x"FF",
	x"00", x"01", x"FF", x"01", x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE",
	x"00", x"00", x"01", x"00", x"FF", x"00", x"FF", x"FE", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FE", x"01", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FE", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"01", x"FF", x"FF", x"00", x"FF", x"FF", x"01",
	x"FF", x"FF", x"FE", x"01", x"FF", x"00", x"FE", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"01", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"00", x"FE",
	x"00", x"FF", x"01", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"FF", x"01",
	x"00", x"01", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FE", x"00", x"00", x"00",
	x"FE", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FE", x"00", x"FE", x"00", x"FF", x"FF", x"00", x"01", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"FF", x"01", x"FF", x"00", x"FE", x"00",
	x"FE", x"00", x"FF", x"01", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"00", x"FE", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"FE", x"00", x"00", x"00", x"00", x"00", x"FE", x"01", x"00", x"00",
	x"FF", x"00", x"FE", x"00", x"FF", x"00", x"FF", x"01", x"FF", x"00", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"01", x"FE",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"01", x"00", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"01", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"01", x"FF", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"01", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"01", x"00", x"FF", x"FF", x"00", x"FF",
	x"01", x"FF", x"FF", x"00", x"01", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"FF", x"01", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"00", x"FF", x"01", x"FF", x"01", x"FE", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"01", x"00", x"FF", x"00", x"FE", x"FF", x"01", x"FF", x"FE", x"01", x"00",
	x"01", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"FF", x"00",
	x"FE", x"00", x"FE", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"01", x"FF", x"FF", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"01", x"FF", x"00", x"00", x"FF", x"FE",
	x"01", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"01",
	x"FF", x"FF", x"FF", x"01", x"FF", x"00", x"FF", x"FF", x"01", x"FF", x"00", x"00",
	x"FF", x"00", x"FF", x"01", x"FE", x"00", x"00", x"01", x"FE", x"00", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"01", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FE", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"FF", x"FE", x"01", x"FF", x"00", x"00", x"FF", x"01", x"00", x"00", x"00",
	x"FE", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"01", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"01", x"FE", x"01", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"FE", x"00", x"FF", x"01", x"FF", x"FF", x"FE", x"01", x"FF", x"FF", x"FF",
	x"01", x"FF", x"01", x"FF", x"FE", x"01", x"FF", x"01", x"FE", x"02", x"FF", x"00",
	x"FF", x"FF", x"FF", x"00", x"01", x"FF", x"FF", x"01", x"01", x"FF", x"00", x"FF",
	x"FF", x"FF", x"01", x"FE", x"00", x"00", x"01", x"FE", x"00", x"00", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"01", x"FF", x"00", x"00", x"FF",
	x"00", x"FF", x"01", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"01", x"FF", x"FE", x"00", x"FF", x"01", x"FD", x"00", x"FF", x"01", x"FE", x"00",
	x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"01", x"FF", x"01", x"FE", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"01", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FE", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FE", x"01", x"FE", x"00", x"FE", x"00",
	x"FE", x"00", x"FE", x"01", x"FE", x"00", x"01", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FE", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"01", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"01", x"FF", x"00", x"FF", x"FF", x"01", x"FE",
	x"00", x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"FE", x"00",
	x"00", x"01", x"FE", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"01", x"00", x"FF", x"00", x"00", x"01", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"01", x"FF", x"00", x"FE", x"00", x"FF", x"01", x"FE", x"01", x"FE",
	x"01", x"FE", x"01", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FE", x"01",
	x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"01", x"FF",
	x"00", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"00", x"00", x"FE", x"01", x"FF",
	x"00", x"00", x"FF", x"00", x"FE", x"00", x"00", x"01", x"FE", x"FF", x"00", x"FE",
	x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"01", x"FE", x"01", x"FF", x"FF", x"00",
	x"FF", x"FF", x"00", x"00", x"FF", x"01", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FE", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"FF",
	x"00", x"FE", x"01", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"01", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"01", x"01",
	x"FF", x"00", x"FE", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FE",
	x"00", x"00", x"FF", x"00", x"FE", x"01", x"FF", x"00", x"FF", x"FF", x"00", x"FF",
	x"FF", x"01", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"01", x"FE", x"01", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"00", x"FE", x"00", x"FF",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"FF", x"01", x"FF", x"01", x"FF", x"00", x"FE", x"FF",
	x"FF", x"01", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"00", x"FF", x"FE", x"01", x"FE", x"00", x"00", x"00", x"FF", x"FF", x"00", x"01",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"FF", x"00", x"FF",
	x"FF", x"FF", x"01", x"00", x"FF", x"00", x"FF", x"01", x"FF", x"00", x"FE", x"00",
	x"FF", x"00", x"00", x"FF", x"01", x"FF", x"00", x"00", x"FE", x"01", x"00", x"FF",
	x"01", x"FE", x"00", x"00", x"00", x"FF", x"FE", x"00", x"01", x"FF", x"00", x"FF",
	x"00", x"FE", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"FF", x"01", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FE", x"00",
	x"00", x"00", x"00", x"FF", x"01", x"FF", x"00", x"FE", x"00", x"FF", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"01", x"FF", x"FE", x"01", x"FF", x"FF", x"FF", x"FE",
	x"00", x"FF", x"01", x"FF", x"FF", x"FF", x"FF", x"00", x"FE", x"FF", x"00", x"00",
	x"00", x"00", x"FE", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"01", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FE", x"01", x"FF", x"00", x"FF",
	x"FF", x"FE", x"00", x"FF", x"FF", x"00", x"FF", x"01", x"FE", x"00", x"FE", x"00",
	x"FF", x"00", x"FF", x"01", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"01", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF",
	x"FF", x"01", x"00", x"00", x"01", x"FF", x"01", x"FE", x"01", x"FE", x"00", x"FF",
	x"00", x"FF", x"FF", x"01", x"00", x"FF", x"00", x"FF", x"FF", x"01", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FE",
	x"00", x"00", x"FF", x"01", x"FF", x"00", x"01", x"FF", x"00", x"FE", x"00", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"FE", x"00", x"FF", x"00", x"FE", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FE",
	x"01", x"FF", x"00", x"FE", x"FF", x"00", x"FF", x"01", x"FF", x"00", x"FF", x"FF",
	x"FE", x"00", x"FF", x"00", x"00", x"00", x"FE", x"00", x"FE", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"01", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FE", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FE", x"FF",
	x"00", x"01", x"FF", x"00", x"FE", x"00", x"FF", x"00", x"FE", x"FF", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FE", x"01", x"FE", x"00", x"01", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FE", x"00", x"FF", x"01", x"FE", x"00", x"FF", x"00", x"FF", x"01", x"FF", x"FF",
	x"01", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"01", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FE", x"01", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FE", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"01", x"FE", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"01", x"FF", x"00", x"00", x"FE", x"01", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"01", x"FF",
	x"01", x"FF", x"00", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF",
	x"01", x"00", x"FE", x"01", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"01", x"FF",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FE", x"00", x"FF", x"00", x"FF", x"00", x"01", x"FF", x"FF", x"FE", x"00", x"FF",
	x"FF", x"01", x"FF", x"FF", x"00", x"00", x"FE", x"00", x"FE", x"00", x"00", x"01",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"00", x"FE", x"00", x"00", x"FF", x"01", x"FE", x"00", x"FF", x"FF", x"01",
	x"FF", x"FF", x"01", x"FF", x"00", x"FF", x"01", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FE", x"FF", x"00", x"FF", x"00", x"FE", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"FE", x"00", x"FF", x"01", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"01", x"FE", x"00", x"00", x"00", x"FF", x"00", x"FF", x"01",
	x"00", x"FF", x"FF", x"00", x"01", x"FF", x"00", x"FE", x"00", x"FF", x"FF", x"FE",
	x"00", x"00", x"01", x"FE", x"00", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"01",
	x"FE", x"01", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"01", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE",
	x"00", x"FE", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"01", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"FF", x"00", x"FF", x"01", x"00", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"00", x"FF", x"01", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FE", x"00", x"00", x"FF", x"01", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"FF",
	x"01", x"FF", x"00", x"00", x"FE", x"00", x"FF", x"00", x"00", x"00", x"01", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FE", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"FE", x"FF", x"00", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"FF", x"01", x"FF", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FF", x"00",
	x"FF", x"FE", x"01", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"01", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FE", x"00", x"FF", x"01", x"FF",
	x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"FE", x"01",
	x"FE", x"00", x"FE", x"00", x"FF", x"00", x"FE", x"00", x"FE", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"FE", x"01", x"FF", x"00", x"FE", x"00",
	x"00", x"FF", x"FF", x"FF", x"01", x"FF", x"00", x"00", x"FE", x"01", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"FF",
	x"01", x"00", x"00", x"FE", x"00", x"FF", x"00", x"00", x"00", x"FE", x"00", x"FF",
	x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"00", x"01", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FE", x"01", x"FE", x"00", x"FE", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FE", x"01", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FE", x"00", x"FF",
	x"00", x"00", x"FE", x"FF", x"00", x"00", x"00", x"FE", x"00", x"FF", x"00", x"FE",
	x"FF", x"FF", x"FF", x"00", x"00", x"FE", x"01", x"FE", x"01", x"FE", x"00", x"00",
	x"FF", x"FF", x"00", x"FF", x"01", x"00", x"FF", x"00", x"FE", x"00", x"FE", x"00",
	x"00", x"FF", x"01", x"FF", x"00", x"FE", x"01", x"FE", x"00", x"00", x"FE", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"FE", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"FF", x"01", x"FF", x"00", x"FF", x"FF", x"01", x"FF", x"01", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"01", x"FF", x"00", x"00", x"FE", x"00", x"00",
	x"FE", x"00", x"FE", x"00", x"FF", x"00", x"FE", x"00", x"FF", x"01", x"FE", x"00",
	x"FF", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"FF", x"01", x"00", x"00", x"FF", x"01", x"FE", x"00", x"FF", x"FF",
	x"01", x"FF", x"00", x"FF", x"FF", x"01", x"FE", x"00", x"FF", x"00", x"FF", x"FF",
	x"01", x"FF", x"FF", x"01", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF",
	x"FF", x"00", x"00", x"FF", x"00", x"FF", x"01", x"FE", x"00", x"00", x"FF", x"01",
	x"FE", x"00", x"FF", x"00", x"FF", x"FF", x"01", x"FF", x"FF", x"01", x"FE", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"FE", x"00", x"00", x"FF", x"00", x"FE", x"01", x"FE", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"FF", x"00", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00",
	x"FE", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FE", x"FF", x"00", x"FE", x"00",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FE", x"00", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"01", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"01", x"00", x"01", x"FE",
	x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"01", x"FE", x"01", x"00", x"00", x"00", x"FE", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"FF", x"00", x"FE", x"01", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"FE", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FE",
	x"00", x"FF", x"01", x"FF", x"00", x"00", x"FE", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"01", x"FE", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FE", x"00", x"00", x"FE", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"01", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FE", x"01",
	x"FF", x"FF", x"00", x"00", x"00", x"FE", x"00", x"FF", x"00", x"00", x"00", x"FF",
	x"00", x"FE", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF",
	x"01", x"FE", x"FF", x"FF", x"FF", x"01", x"FF", x"01", x"FE", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"FE", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"FF", x"01", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF",
	x"01", x"FF", x"00", x"FE", x"00", x"00", x"FF", x"FF", x"FE", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FE",
	x"00", x"FF", x"FF", x"01", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"01", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FE", x"00", x"FF", x"00", x"FF", x"FF",
	x"FE", x"01", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"00", x"01", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"01", x"FF",
	x"00", x"FF", x"00", x"01", x"FF", x"00", x"00", x"FE", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"FE", x"FF", x"00", x"01", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"FE", x"00", x"FF", x"01", x"00", x"FF", x"01", x"FE", x"01", x"00", x"FE", x"01",
	x"00", x"FF", x"00", x"FF", x"00", x"FE", x"01", x"FF", x"01", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"01",
	x"FF", x"FE", x"00", x"FF", x"00", x"01", x"FF", x"FE", x"00", x"01", x"FF", x"FF",
	x"FE", x"00", x"FF", x"00", x"00", x"FE", x"00", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"FF", x"00", x"FE", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"01", x"FF", x"00",
	x"FE", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"00", x"01", x"FF", x"FF",
	x"01", x"FE", x"00", x"FF", x"FF", x"01", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"01", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"00", x"FF", x"00",
	x"FE", x"00", x"FF", x"01", x"00", x"FF", x"00", x"FE", x"00", x"00", x"FF", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"01", x"FF", x"00", x"FF", x"00", x"FE", x"00", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"01", x"FF", x"00", x"FF", x"FF", x"00", x"01", x"00", x"00", x"FE", x"01", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FE", x"00", x"FF", x"00", x"FF",
	x"00", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"01", x"00", x"00", x"00", x"FE",
	x"01", x"FF", x"01", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"01", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"00", x"FF", x"01",
	x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"01", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"FE", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF"
	);
	
signal cnt_out: unsigned(15 downto 0) := (others => '0');	
signal play_sound: std_logic := '0';
constant cnt_max: integer := 18687;
signal out_signal: signed(7 downto 0) := x"00";

begin
	
process (CLK)
begin
    if rising_edge(CLK) then
        if RST = '1' then
            play_sound <= '0';
        elsif PLAY = '1' then
            play_sound <= '1';
        elsif PLAY = '0' and cnt_out = cnt_max then
            play_sound <= '0';
        end if;
    end if;
end process;

	
-- 12bit counter
process (CLK)
begin     
    if rising_edge(CLK) then
        if RST = '1' then
            cnt_out <= (others => '0');
        elsif CE = '1' and play_sound = '1' then
            cnt_out <= cnt_out + 1;       
        end if;
        if cnt_out = cnt_max then
            cnt_out <= (others => '0');            
        end if;        
    end if;
end process;

process (CLK) 
begin
    if rising_edge(CLK) then
        if RST = '1' then
            out_signal <= x"00";
        elsif CE = '1' then
            out_signal <= crash_sound(conv_integer(cnt_out));
        end if;
    end if;    
end process;

SAMPLE_OUT <= out_signal;

end Behavioral;




