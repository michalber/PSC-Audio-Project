----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 25.12.2018 17:39:59
-- Design Name: 
-- Module Name: Snare - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_1164.ALL;


-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Snare is
    Port ( CLK : in STD_LOGIC;
           CE : in STD_LOGIC;
           RST : in STD_LOGIC;
           PLAY : in STD_LOGIC;
           SNARE_SAMP_O : out signed(7 downto 0)
           );
end Snare;

architecture Behavioral of Snare is

type memory is array (0 to 19212) of signed(7 downto 0);
constant snare_sound: memory := (	
	x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"03", x"04", x"06", x"06", x"01", x"FC",
	x"FB", x"FD", x"00", x"04", x"0A", x"10", x"15", x"19", x"1E", x"23", x"27", x"2A",
	x"2B", x"2B", x"29", x"27", x"26", x"25", x"23", x"22", x"20", x"1F", x"1D", x"1B",
	x"19", x"17", x"15", x"13", x"13", x"14", x"10", x"0A", x"06", x"FE", x"F7", x"EF",
	x"E9", x"F5", x"0E", x"22", x"21", x"05", x"E5", x"D1", x"C5", x"BF", x"C0", x"C0",
	x"C1", x"C2", x"C2", x"C2", x"C1", x"BF", x"BF", x"BF", x"C0", x"C2", x"C6", x"C9",
	x"CB", x"CD", x"CE", x"D1", x"D4", x"D9", x"DE", x"E5", x"EC", x"F4", x"FC", x"03",
	x"0A", x"0F", x"13", x"16", x"18", x"19", x"1A", x"1D", x"20", x"22", x"22", x"1D",
	x"17", x"10", x"0B", x"12", x"23", x"27", x"20", x"1A", x"12", x"07", x"FB", x"F6",
	x"F9", x"FB", x"FB", x"F8", x"F2", x"E7", x"DB", x"D5", x"D5", x"DB", x"DE", x"DE",
	x"D7", x"C9", x"C8", x"CA", x"D1", x"F9", x"2A", x"40", x"3F", x"3B", x"33", x"30",
	x"29", x"10", x"0D", x"01", x"F3", x"F8", x"EA", x"EA", x"F7", x"0D", x"36", x"56",
	x"63", x"5F", x"5A", x"47", x"2C", x"1E", x"1A", x"2B", x"3D", x"4E", x"60", x"6C",
	x"76", x"76", x"74", x"73", x"71", x"6F", x"6D", x"6D", x"6B", x"69", x"66", x"59",
	x"3E", x"23", x"0C", x"F9", x"ED", x"E3", x"E0", x"DF", x"E1", x"E5", x"E2", x"D9",
	x"D1", x"D3", x"D8", x"E7", x"F6", x"FD", x"FF", x"00", x"06", x"0A", x"07", x"05",
	x"01", x"00", x"FF", x"FF", x"FE", x"F1", x"D6", x"BF", x"BC", x"C4", x"CD", x"D6",
	x"E5", x"F9", x"0D", x"1E", x"2A", x"32", x"36", x"39", x"39", x"38", x"35", x"32",
	x"2E", x"2B", x"27", x"21", x"1C", x"19", x"17", x"14", x"11", x"0D", x"08", x"02",
	x"FF", x"00", x"02", x"05", x"05", x"FF", x"F5", x"E6", x"D4", x"C2", x"B5", x"AE",
	x"B5", x"C8", x"D5", x"D9", x"D6", x"CB", x"B9", x"A5", x"9B", x"9C", x"9F", x"A1",
	x"A3", x"A6", x"A8", x"AA", x"AB", x"AA", x"A8", x"AF", x"C0", x"D5", x"E4", x"F1",
	x"FF", x"10", x"26", x"37", x"37", x"29", x"17", x"02", x"ED", x"D9", x"CB", x"C5",
	x"C6", x"C9", x"CD", x"D4", x"DD", x"EB", x"F3", x"FA", x"05", x"F2", x"E1", x"E8",
	x"F0", x"1C", x"52", x"5D", x"53", x"45", x"38", x"2D", x"1E", x"12", x"08", x"03",
	x"FF", x"00", x"F4", x"E1", x"DC", x"DD", x"F8", x"14", x"25", x"30", x"2B", x"24",
	x"19", x"13", x"11", x"12", x"1B", x"26", x"2F", x"2B", x"2C", x"2A", x"29", x"35",
	x"3B", x"39", x"2D", x"28", x"2A", x"29", x"2A", x"2C", x"35", x"3A", x"41", x"48",
	x"4D", x"51", x"4F", x"50", x"50", x"4C", x"3F", x"2D", x"1F", x"10", x"05", x"FE",
	x"FE", x"07", x"1B", x"36", x"45", x"47", x"40", x"35", x"2A", x"23", x"20", x"26",
	x"31", x"3D", x"48", x"51", x"5E", x"6C", x"72", x"73", x"73", x"69", x"56", x"45",
	x"3C", x"3D", x"41", x"45", x"4A", x"4E", x"51", x"53", x"55", x"56", x"55", x"52",
	x"4E", x"49", x"3F", x"33", x"27", x"1C", x"1C", x"2A", x"3A", x"40", x"36", x"1D",
	x"FF", x"DF", x"C0", x"AA", x"A6", x"A9", x"AB", x"B3", x"C0", x"CD", x"D5", x"D5",
	x"D0", x"C5", x"B9", x"B0", x"AF", x"AF", x"AF", x"B0", x"B8", x"CA", x"E0", x"FA",
	x"17", x"31", x"4A", x"59", x"5E", x"5C", x"56", x"4D", x"44", x"3D", x"3B", x"39",
	x"35", x"2F", x"26", x"1C", x"13", x"0B", x"07", x"05", x"05", x"06", x"03", x"FD",
	x"F4", x"E9", x"DD", x"D4", x"CC", x"C4", x"C1", x"C4", x"C5", x"C1", x"BE", x"BD",
	x"B9", x"B1", x"A6", x"99", x"92", x"91", x"92", x"92", x"91", x"8F", x"8D", x"8E",
	x"93", x"97", x"9B", x"9F", x"A3", x"A5", x"A7", x"AA", x"AD", x"B0", x"B2", x"B5",
	x"B8", x"BB", x"C0", x"C5", x"CB", x"CF", x"D2", x"D3", x"D5", x"DA", x"E4", x"F2",
	x"00", x"0E", x"18", x"0D", x"FE", x"06", x"13", x"15", x"1D", x"25", x"28", x"27",
	x"24", x"24", x"23", x"20", x"1D", x"1A", x"18", x"19", x"1B", x"1C", x"19", x"16",
	x"15", x"15", x"18", x"1D", x"1B", x"05", x"FA", x"E5", x"B9", x"CA", x"EB", x"F3",
	x"DA", x"B8", x"DD", x"FD", x"FD", x"01", x"FD", x"FD", x"FC", x"FF", x"F9", x"F5",
	x"E6", x"C8", x"B7", x"C3", x"EF", x"05", x"18", x"37", x"3F", x"46", x"4F", x"5B",
	x"5E", x"5B", x"5F", x"63", x"66", x"60", x"5C", x"5E", x"5E", x"59", x"5A", x"61",
	x"62", x"62", x"60", x"56", x"48", x"42", x"3C", x"38", x"3E", x"43", x"41", x"3C",
	x"3F", x"46", x"45", x"3E", x"3E", x"3D", x"2D", x"20", x"20", x"26", x"28", x"1F",
	x"18", x"15", x"10", x"07", x"05", x"0F", x"16", x"19", x"1A", x"1B", x"1A", x"0D",
	x"08", x"0E", x"03", x"EE", x"E4", x"E4", x"E6", x"E8", x"EB", x"E9", x"E7", x"E4",
	x"D6", x"CB", x"C4", x"C0", x"C1", x"C5", x"CF", x"E2", x"EB", x"E0", x"CB", x"BC",
	x"AE", x"A3", x"A1", x"A0", x"A2", x"AA", x"B6", x"C2", x"C3", x"B5", x"A7", x"A9",
	x"B3", x"B1", x"B1", x"BF", x"D2", x"E1", x"ED", x"F1", x"F5", x"FD", x"04", x"10",
	x"1C", x"15", x"05", x"F8", x"F2", x"F6", x"FB", x"02", x"0B", x"12", x"16", x"17",
	x"13", x"10", x"1E", x"36", x"4D", x"48", x"27", x"1C", x"1F", x"14", x"04", x"F2",
	x"E0", x"D7", x"D1", x"C3", x"B3", x"AA", x"AB", x"B4", x"B6", x"B4", x"BA", x"C2",
	x"C2", x"BA", x"B4", x"B9", x"C1", x"BB", x"AF", x"B8", x"CD", x"E1", x"EB", x"EB",
	x"F2", x"F6", x"EF", x"F1", x"F6", x"FC", x"08", x"12", x"1F", x"2F", x"39", x"38",
	x"36", x"3C", x"42", x"46", x"45", x"4A", x"5E", x"72", x"71", x"67", x"66", x"6D",
	x"7A", x"7F", x"7F", x"7F", x"7F", x"7B", x"6C", x"55", x"47", x"42", x"3B", x"32",
	x"2B", x"1D", x"03", x"F5", x"1D", x"3F", x"23", x"1F", x"4D", x"5A", x"33", x"10",
	x"0D", x"04", x"0D", x"2C", x"2E", x"28", x"29", x"20", x"03", x"D9", x"CF", x"D2",
	x"BE", x"AB", x"AB", x"B9", x"CF", x"E8", x"FF", x"14", x"25", x"32", x"39", x"3A",
	x"3D", x"43", x"46", x"45", x"44", x"43", x"3B", x"38", x"39", x"3A", x"3B", x"3C",
	x"39", x"39", x"45", x"45", x"3C", x"3B", x"3D", x"3D", x"2F", x"20", x"1A", x"1B",
	x"16", x"0B", x"05", x"05", x"02", x"F4", x"E9", x"E9", x"F1", x"FF", x"F7", x"DD",
	x"CA", x"C3", x"CA", x"CF", x"CD", x"CD", x"D2", x"D0", x"C9", x"CA", x"C3", x"B6",
	x"B3", x"B4", x"B5", x"B4", x"B7", x"C2", x"D2", x"E0", x"ED", x"02", x"12", x"14",
	x"10", x"09", x"06", x"0B", x"10", x"10", x"0E", x"0A", x"04", x"FF", x"FB", x"F6",
	x"F4", x"F5", x"F2", x"F3", x"FC", x"02", x"FB", x"E1", x"D0", x"D2", x"CD", x"C6",
	x"C5", x"B9", x"A7", x"A0", x"A6", x"A9", x"AD", x"B2", x"B3", x"B1", x"AC", x"A8",
	x"AD", x"B0", x"AC", x"A5", x"9F", x"9F", x"AC", x"B8", x"B1", x"A6", x"A5", x"A9",
	x"C0", x"DE", x"F7", x"13", x"29", x"2B", x"1F", x"19", x"25", x"34", x"3A", x"38",
	x"32", x"31", x"31", x"35", x"35", x"32", x"37", x"3E", x"41", x"40", x"3B", x"33",
	x"1F", x"0E", x"09", x"DB", x"AC", x"C8", x"E3", x"EB", x"EC", x"E1", x"EC", x"ED",
	x"F4", x"FC", x"EE", x"E5", x"E0", x"E3", x"DE", x"EC", x"01", x"08", x"0E", x"0A",
	x"13", x"19", x"25", x"37", x"3E", x"45", x"4A", x"55", x"56", x"56", x"57", x"54",
	x"55", x"54", x"54", x"4D", x"45", x"3D", x"2E", x"2D", x"30", x"36", x"3A", x"48",
	x"5D", x"6E", x"78", x"73", x"6F", x"71", x"72", x"73", x"74", x"79", x"77", x"6C",
	x"55", x"3D", x"2C", x"1C", x"18", x"1B", x"18", x"11", x"08", x"05", x"0A", x"16",
	x"18", x"04", x"F3", x"F9", x"FC", x"F8", x"F3", x"EB", x"F6", x"08", x"0B", x"0C",
	x"0A", x"04", x"06", x"0C", x"0D", x"12", x"1F", x"1D", x"13", x"18", x"27", x"30",
	x"3E", x"4B", x"51", x"4F", x"49", x"48", x"48", x"46", x"45", x"49", x"45", x"35",
	x"2C", x"24", x"1C", x"19", x"16", x"15", x"10", x"09", x"03", x"00", x"0A", x"1A",
	x"1A", x"0F", x"10", x"0E", x"F5", x"DF", x"E2", x"E4", x"D7", x"D2", x"D9", x"DE",
	x"D5", x"C9", x"C6", x"C5", x"CC", x"D9", x"E6", x"F0", x"EC", x"DC", x"C5", x"B4",
	x"B7", x"BF", x"B7", x"B0", x"B3", x"B9", x"BE", x"C2", x"D6", x"FF", x"19", x"12",
	x"0B", x"09", x"F7", x"E2", x"E8", x"04", x"09", x"FB", x"F6", x"EA", x"E8", x"F4",
	x"F9", x"02", x"13", x"1E", x"18", x"08", x"02", x"F7", x"E3", x"D3", x"C9", x"BE",
	x"B6", x"B3", x"BB", x"CB", x"D2", x"CA", x"BC", x"C2", x"DD", x"F1", x"F6", x"FE",
	x"13", x"20", x"1A", x"08", x"EE", x"D3", x"BC", x"AE", x"A8", x"A9", x"B0", x"BA",
	x"BD", x"B5", x"B0", x"AC", x"AE", x"C1", x"DB", x"F0", x"F4", x"EF", x"FA", x"07",
	x"11", x"1D", x"28", x"31", x"2D", x"21", x"19", x"10", x"09", x"0A", x"08", x"F7",
	x"EA", x"E9", x"E7", x"E4", x"DC", x"D1", x"D3", x"CA", x"BC", x"BD", x"C7", x"D1",
	x"D1", x"D6", x"E6", x"FC", x"13", x"1B", x"19", x"17", x"12", x"0C", x"07", x"07",
	x"05", x"FE", x"FB", x"04", x"11", x"20", x"2F", x"28", x"19", x"1B", x"23", x"24",
	x"21", x"27", x"32", x"44", x"63", x"78", x"7D", x"7B", x"74", x"6E", x"6F", x"72",
	x"70", x"67", x"66", x"6B", x"6F", x"78", x"78", x"63", x"46", x"3B", x"4B", x"50",
	x"3B", x"2E", x"3A", x"4A", x"48", x"39", x"2D", x"28", x"1E", x"0C", x"F8", x"EB",
	x"EA", x"E9", x"DD", x"D4", x"E0", x"EE", x"ED", x"EC", x"EC", x"E7", x"E7", x"ED",
	x"F7", x"02", x"0A", x"0C", x"0C", x"0C", x"0E", x"10", x"0C", x"0D", x"16", x"1B",
	x"15", x"0A", x"02", x"02", x"09", x"10", x"1B", x"23", x"1C", x"10", x"06", x"0B",
	x"1C", x"1E", x"0C", x"F5", x"E5", x"E1", x"E7", x"F6", x"F9", x"F3", x"EE", x"DD",
	x"C9", x"C7", x"D2", x"DA", x"DF", x"DC", x"D3", x"CA", x"C2", x"BC", x"B5", x"AB",
	x"A8", x"A7", x"A3", x"A7", x"B2", x"BF", x"CE", x"D5", x"D9", x"E0", x"E7", x"E8",
	x"DB", x"C8", x"BD", x"C1", x"D2", x"E4", x"F2", x"F9", x"00", x"01", x"FB", x"F6",
	x"F0", x"E8", x"E6", x"E6", x"E3", x"E9", x"FA", x"0F", x"1E", x"27", x"2B", x"2F",
	x"34", x"33", x"34", x"37", x"2D", x"1B", x"13", x"17", x"06", x"E8", x"E5", x"F3",
	x"FB", x"F7", x"E6", x"D5", x"CD", x"C9", x"C5", x"C0", x"C4", x"CB", x"C4", x"BD",
	x"BA", x"B1", x"AD", x"BC", x"CC", x"CA", x"C2", x"B3", x"AA", x"B9", x"D1", x"DC",
	x"D6", x"D3", x"D2", x"C9", x"C0", x"C5", x"DA", x"F5", x"09", x"03", x"F8", x"F8",
	x"FA", x"F5", x"F5", x"01", x"03", x"00", x"09", x"0F", x"16", x"28", x"3F", x"50",
	x"53", x"4C", x"44", x"34", x"1C", x"10", x"08", x"F5", x"E6", x"EF", x"FE", x"00",
	x"04", x"13", x"1F", x"1E", x"1F", x"27", x"2F", x"33", x"2F", x"2B", x"2D", x"33",
	x"36", x"30", x"27", x"24", x"26", x"25", x"1A", x"09", x"04", x"0E", x"19", x"19",
	x"13", x"1C", x"2D", x"36", x"35", x"25", x"19", x"26", x"3A", x"3B", x"33", x"38",
	x"44", x"4D", x"4B", x"45", x"4A", x"55", x"56", x"4E", x"44", x"39", x"36", x"3A",
	x"39", x"38", x"32", x"25", x"12", x"00", x"F4", x"E9", x"DC", x"CD", x"CC", x"CC",
	x"C5", x"C6", x"C6", x"CA", x"CE", x"DD", x"F0", x"EE", x"EA", x"F1", x"F9", x"F2",
	x"EE", x"F9", x"FA", x"F3", x"F6", x"08", x"1A", x"19", x"0C", x"09", x"13", x"19",
	x"1B", x"19", x"11", x"0C", x"0C", x"0F", x"0F", x"13", x"18", x"16", x"11", x"16",
	x"1D", x"15", x"0C", x"0D", x"08", x"F9", x"E9", x"E5", x"DF", x"D4", x"D1", x"D2",
	x"C9", x"BD", x"BF", x"CB", x"CF", x"C9", x"C3", x"C0", x"B9", x"B5", x"B5", x"B3",
	x"B5", x"BA", x"B0", x"A0", x"9E", x"AC", x"B8", x"C2", x"CE", x"D7", x"D9", x"DB",
	x"DC", x"D8", x"DC", x"DF", x"D8", x"D8", x"E3", x"F2", x"F9", x"F8", x"FF", x"10",
	x"14", x"0E", x"12", x"1C", x"23", x"2A", x"35", x"3B", x"3E", x"37", x"26", x"1F",
	x"21", x"25", x"23", x"17", x"11", x"14", x"1C", x"1E", x"15", x"07", x"F9", x"EE",
	x"E3", x"DC", x"D4", x"CB", x"CA", x"CE", x"D1", x"C7", x"BE", x"CB", x"D9", x"D5",
	x"CF", x"CD", x"D9", x"EC", x"EF", x"E7", x"E3", x"E2", x"DF", x"D3", x"CC", x"D5",
	x"DD", x"D5", x"D3", x"E3", x"EE", x"F2", x"FC", x"05", x"0E", x"15", x"16", x"15",
	x"15", x"1D", x"25", x"29", x"2E", x"34", x"3B", x"3C", x"3B", x"3B", x"31", x"21",
	x"15", x"0B", x"FC", x"FB", x"0B", x"14", x"13", x"07", x"02", x"06", x"01", x"F9",
	x"FE", x"10", x"18", x"0D", x"08", x"13", x"15", x"07", x"FD", x"03", x"0B", x"00",
	x"F3", x"FE", x"10", x"0A", x"F6", x"EC", x"F1", x"F7", x"F2", x"EB", x"EA", x"F0",
	x"FA", x"07", x"1B", x"29", x"21", x"0D", x"FD", x"F3", x"F9", x"0B", x"0D", x"06",
	x"0B", x"18", x"26", x"2B", x"31", x"3A", x"3B", x"37", x"2F", x"29", x"2A", x"2B",
	x"1E", x"0A", x"07", x"0B", x"0C", x"0B", x"0A", x"0A", x"06", x"05", x"05", x"03",
	x"03", x"02", x"00", x"00", x"04", x"0F", x"15", x"0D", x"08", x"13", x"19", x"12",
	x"07", x"01", x"F9", x"ED", x"EE", x"FD", x"0C", x"14", x"0F", x"08", x"07", x"0E",
	x"14", x"0F", x"0B", x"0F", x"16", x"20", x"26", x"22", x"19", x"19", x"1C", x"1A",
	x"12", x"0B", x"0A", x"02", x"F8", x"F4", x"E9", x"D8", x"DB", x"ED", x"F0", x"EB",
	x"EC", x"E8", x"DC", x"D5", x"DD", x"EA", x"F0", x"E9", x"DD", x"DE", x"E4", x"DB",
	x"D3", x"D6", x"E1", x"E8", x"DC", x"CB", x"CA", x"CD", x"CE", x"D2", x"D9", x"DB",
	x"D7", x"D6", x"D5", x"D9", x"DD", x"DA", x"DB", x"E7", x"F4", x"F8", x"04", x"12",
	x"15", x"1A", x"15", x"00", x"F3", x"F7", x"00", x"03", x"0C", x"1E", x"27", x"1F",
	x"18", x"14", x"09", x"F8", x"ED", x"F7", x"03", x"02", x"FC", x"F9", x"F6", x"F0",
	x"EF", x"ED", x"E2", x"DF", x"ED", x"F9", x"EC", x"D5", x"D1", x"D9", x"DA", x"CF",
	x"BD", x"B2", x"B5", x"C7", x"DD", x"E3", x"DF", x"E2", x"EC", x"E9", x"E1", x"E3",
	x"E9", x"EB", x"E4", x"DF", x"E2", x"EB", x"00", x"15", x"1A", x"0D", x"06", x"14",
	x"22", x"22", x"1E", x"23", x"2C", x"31", x"2F", x"2F", x"33", x"2D", x"21", x"21",
	x"25", x"20", x"17", x"18", x"17", x"11", x"0F", x"11", x"16", x"1D", x"1B", x"14",
	x"10", x"0F", x"0E", x"0A", x"08", x"03", x"F5", x"EE", x"EF", x"ED", x"EC", x"F2",
	x"F7", x"F9", x"F9", x"F5", x"EE", x"ED", x"EE", x"ED", x"EB", x"E8", x"E2", x"E0",
	x"E3", x"EB", x"F1", x"F0", x"F0", x"F8", x"FF", x"FB", x"EE", x"EA", x"FB", x"0F",
	x"17", x"1E", x"29", x"37", x"41", x"44", x"45", x"47", x"42", x"39", x"37", x"39",
	x"32", x"28", x"26", x"28", x"29", x"2A", x"2E", x"30", x"22", x"12", x"15", x"1D",
	x"15", x"03", x"FA", x"F5", x"F6", x"FE", x"04", x"09", x"0F", x"12", x"0A", x"FB",
	x"F9", x"FE", x"02", x"06", x"09", x"0A", x"0E", x"11", x"13", x"11", x"0C", x"0A",
	x"03", x"FA", x"F7", x"F9", x"F7", x"F0", x"EA", x"E2", x"E0", x"E6", x"E5", x"DC",
	x"D8", x"E1", x"EB", x"EF", x"F4", x"F9", x"F7", x"EE", x"F2", x"FD", x"FC", x"F8",
	x"FF", x"04", x"F6", x"DD", x"D2", x"DE", x"F0", x"F9", x"F7", x"F8", x"01", x"01",
	x"FA", x"F2", x"EF", x"F0", x"EA", x"E1", x"E5", x"EC", x"EC", x"E6", x"DE", x"DC",
	x"DE", x"E7", x"F5", x"F0", x"E2", x"E2", x"EF", x"F5", x"F2", x"F7", x"FD", x"FE",
	x"FB", x"FD", x"01", x"FB", x"F4", x"FB", x"09", x"0A", x"00", x"02", x"11", x"1C",
	x"1E", x"1A", x"1B", x"24", x"1F", x"10", x"0F", x"11", x"09", x"F4", x"E3", x"E7",
	x"F3", x"F1", x"E8", x"E0", x"D9", x"D3", x"D4", x"D8", x"DC", x"E1", x"E0", x"D7",
	x"CE", x"CC", x"D1", x"D7", x"E3", x"F0", x"F5", x"F5", x"F2", x"F7", x"01", x"04",
	x"06", x"0A", x"0F", x"17", x"13", x"0C", x"15", x"18", x"06", x"F8", x"FF", x"0C",
	x"0D", x"05", x"02", x"00", x"01", x"03", x"FF", x"03", x"10", x"15", x"0B", x"03",
	x"02", x"FB", x"F8", x"04", x"08", x"FD", x"F4", x"F6", x"FB", x"FE", x"FE", x"02",
	x"03", x"FB", x"F6", x"FA", x"00", x"05", x"08", x"05", x"FD", x"00", x"12", x"25",
	x"23", x"1A", x"20", x"30", x"3C", x"31", x"17", x"0D", x"15", x"16", x"09", x"FA",
	x"F9", x"FF", x"F7", x"EF", x"F4", x"F8", x"ED", x"E1", x"E3", x"F0", x"FB", x"01",
	x"04", x"0A", x"11", x"13", x"11", x"16", x"26", x"33", x"38", x"3E", x"3D", x"3B",
	x"45", x"50", x"4E", x"42", x"31", x"22", x"26", x"33", x"34", x"25", x"14", x"0F",
	x"10", x"0F", x"10", x"18", x"21", x"24", x"26", x"22", x"13", x"03", x"FC", x"F8",
	x"F2", x"EE", x"F2", x"03", x"1C", x"24", x"24", x"29", x"29", x"1B", x"0A", x"07",
	x"09", x"FC", x"EA", x"E7", x"F3", x"FC", x"F6", x"EC", x"E8", x"EB", x"ED", x"EA",
	x"E9", x"EA", x"EB", x"EC", x"EB", x"EF", x"F2", x"EA", x"E3", x"EA", x"F5", x"F7",
	x"EE", x"E3", x"DD", x"DD", x"DF", x"E2", x"E7", x"EF", x"FA", x"FA", x"E9", x"E2",
	x"EA", x"F1", x"EE", x"EB", x"EE", x"ED", x"EE", x"FB", x"0A", x"0C", x"06", x"02",
	x"FE", x"F4", x"EA", x"E9", x"EE", x"EE", x"E4", x"E2", x"F3", x"04", x"07", x"FC",
	x"EF", x"EA", x"EC", x"E8", x"D9", x"C9", x"C7", x"CF", x"D7", x"D9", x"D8", x"DD",
	x"EA", x"F0", x"EA", x"E7", x"E8", x"E6", x"DD", x"D4", x"D6", x"E2", x"ED", x"EF",
	x"E8", x"E7", x"F1", x"FE", x"06", x"04", x"03", x"09", x"0B", x"0D", x"0F", x"05",
	x"F7", x"EF", x"EF", x"EF", x"E8", x"E9", x"ED", x"F4", x"F8", x"EB", x"E0", x"E0",
	x"DE", x"D9", x"DC", x"EF", x"05", x"0C", x"0A", x"16", x"28", x"2C", x"24", x"1C",
	x"21", x"2B", x"28", x"1E", x"1F", x"24", x"20", x"1C", x"22", x"2A", x"20", x"0E",
	x"10", x"1B", x"19", x"0A", x"01", x"07", x"14", x"18", x"0E", x"0F", x"17", x"17",
	x"14", x"14", x"17", x"14", x"0C", x"0D", x"19", x"1F", x"18", x"0D", x"07", x"09",
	x"05", x"FA", x"FB", x"08", x"0E", x"0A", x"0A", x"0D", x"11", x"10", x"0F", x"14",
	x"15", x"0F", x"0C", x"13", x"18", x"0F", x"07", x"12", x"27", x"2C", x"25", x"26",
	x"23", x"19", x"11", x"0E", x"11", x"14", x"09", x"FA", x"FA", x"07", x"13", x"16",
	x"14", x"12", x"12", x"10", x"0A", x"06", x"07", x"0C", x"08", x"F9", x"F2", x"F0",
	x"E7", x"E6", x"EE", x"F3", x"ED", x"E5", x"E4", x"E9", x"E8", x"E5", x"EA", x"EE",
	x"EF", x"F4", x"FE", x"05", x"0B", x"12", x"12", x"07", x"F9", x"F5", x"FC", x"FF",
	x"F8", x"EE", x"E6", x"E4", x"E8", x"EB", x"EE", x"EF", x"E8", x"E2", x"E9", x"EB",
	x"E1", x"DA", x"DF", x"E5", x"E6", x"E7", x"EC", x"F4", x"F8", x"F7", x"F5", x"F7",
	x"05", x"10", x"0D", x"06", x"01", x"02", x"02", x"FB", x"F2", x"ED", x"F1", x"F9",
	x"FE", x"FF", x"FD", x"FC", x"F7", x"EC", x"EA", x"F5", x"FC", x"F5", x"F1", x"FD",
	x"0E", x"16", x"12", x"04", x"F7", x"01", x"11", x"0A", x"FB", x"FA", x"FF", x"02",
	x"FE", x"F9", x"FC", x"FD", x"F4", x"EA", x"E3", x"D6", x"CD", x"D2", x"D8", x"D8",
	x"DE", x"EC", x"F6", x"FF", x"01", x"F9", x"EF", x"E2", x"E5", x"FC", x"06", x"00",
	x"F7", x"F8", x"F9", x"F7", x"00", x"03", x"F7", x"F2", x"F2", x"F1", x"ED", x"E9",
	x"EF", x"FB", x"00", x"FC", x"FB", x"FE", x"01", x"02", x"03", x"03", x"FD", x"FC",
	x"05", x"10", x"10", x"0C", x"0F", x"16", x"1B", x"18", x"0F", x"0B", x"0F", x"14",
	x"0F", x"02", x"FA", x"F6", x"F4", x"F6", x"FC", x"0A", x"17", x"18", x"13", x"14",
	x"13", x"08", x"06", x"12", x"19", x"15", x"11", x"14", x"14", x"0C", x"03", x"04",
	x"0A", x"0B", x"08", x"04", x"FF", x"FE", x"FF", x"FE", x"01", x"0F", x"16", x"0E",
	x"0B", x"14", x"1E", x"1B", x"17", x"1B", x"1A", x"13", x"0B", x"02", x"FE", x"01",
	x"02", x"FD", x"F2", x"EF", x"F6", x"FA", x"F5", x"F5", x"01", x"0E", x"0C", x"07",
	x"0F", x"14", x"12", x"11", x"15", x"1B", x"1B", x"19", x"1C", x"16", x"09", x"08",
	x"11", x"17", x"12", x"12", x"1E", x"1E", x"16", x"11", x"08", x"00", x"FF", x"04",
	x"03", x"FE", x"04", x"18", x"25", x"23", x"1A", x"13", x"0D", x"05", x"01", x"02",
	x"02", x"06", x"0D", x"0D", x"0A", x"06", x"FD", x"F7", x"F4", x"F2", x"EF", x"F1",
	x"F4", x"F2", x"EF", x"EC", x"F2", x"00", x"02", x"F5", x"EF", x"F7", x"FC", x"F4",
	x"EC", x"EF", x"F4", x"EE", x"E9", x"F0", x"FF", x"03", x"FD", x"FB", x"00", x"FE",
	x"EF", x"E8", x"EF", x"F2", x"F0", x"EC", x"EA", x"EB", x"ED", x"E7", x"E3", x"EB",
	x"F0", x"E3", x"D6", x"DB", x"E8", x"EA", x"EC", x"F0", x"F1", x"F4", x"F6", x"F4",
	x"F2", x"F3", x"F4", x"F1", x"F1", x"F7", x"F6", x"EF", x"EE", x"F1", x"EC", x"E5",
	x"EC", x"F9", x"03", x"05", x"FF", x"FA", x"F6", x"F2", x"F1", x"F3", x"EE", x"E2",
	x"DA", x"DB", x"DE", x"E1", x"E8", x"ED", x"EC", x"F1", x"FD", x"08", x"0B", x"08",
	x"0D", x"13", x"10", x"10", x"16", x"19", x"12", x"0E", x"12", x"1B", x"1C", x"13",
	x"10", x"13", x"0D", x"05", x"04", x"07", x"0D", x"18", x"21", x"1F", x"11", x"09",
	x"0F", x"13", x"13", x"13", x"11", x"0C", x"07", x"08", x"08", x"FE", x"F6", x"F9",
	x"F9", x"F4", x"F4", x"F8", x"FB", x"FE", x"FE", x"F9", x"EF", x"E7", x"E5", x"ED",
	x"F6", x"FD", x"02", x"FF", x"FC", x"00", x"07", x"08", x"02", x"FB", x"F9", x"FA",
	x"F9", x"F9", x"FF", x"07", x"0B", x"11", x"16", x"12", x"0B", x"08", x"10", x"1A",
	x"16", x"0C", x"0D", x"0F", x"08", x"00", x"FE", x"08", x"0D", x"04", x"00", x"08",
	x"13", x"13", x"0A", x"06", x"09", x"08", x"05", x"0A", x"0D", x"0F", x"14", x"13",
	x"0B", x"07", x"09", x"07", x"02", x"00", x"FD", x"FC", x"FD", x"FE", x"FF", x"03",
	x"07", x"06", x"02", x"05", x"0C", x"11", x"14", x"15", x"0D", x"04", x"02", x"03",
	x"04", x"02", x"FF", x"05", x"0B", x"FE", x"F1", x"EF", x"F3", x"F1", x"E7", x"E4",
	x"E9", x"F0", x"F6", x"F7", x"F6", x"F6", x"F7", x"F8", x"F6", x"F5", x"FA", x"FC",
	x"F4", x"EA", x"E6", x"E3", x"DD", x"DC", x"E6", x"EF", x"EE", x"F2", x"FA", x"FC",
	x"FB", x"F7", x"F5", x"F2", x"EE", x"F3", x"01", x"0A", x"02", x"FB", x"FF", x"05",
	x"06", x"FE", x"F5", x"F4", x"F7", x"F6", x"F3", x"FA", x"02", x"05", x"05", x"02",
	x"FD", x"F8", x"F3", x"F4", x"FC", x"FF", x"F2", x"E4", x"E4", x"EB", x"F0", x"F5",
	x"F9", x"FB", x"04", x"10", x"11", x"09", x"05", x"00", x"F8", x"EA", x"DF", x"EC",
	x"FE", x"FE", x"00", x"04", x"04", x"04", x"0A", x"14", x"15", x"10", x"12", x"16",
	x"12", x"03", x"FE", x"03", x"04", x"FC", x"F4", x"F5", x"FD", x"FF", x"FE", x"04",
	x"05", x"FC", x"F5", x"F6", x"FC", x"04", x"0A", x"0D", x"11", x"0D", x"03", x"FD",
	x"FB", x"F8", x"FB", x"03", x"FC", x"F0", x"F2", x"F8", x"02", x"09", x"0C", x"0D",
	x"09", x"03", x"00", x"01", x"04", x"FF", x"FA", x"00", x"03", x"06", x"0D", x"0F",
	x"0C", x"08", x"08", x"08", x"00", x"F6", x"F4", x"F8", x"F9", x"F4", x"EE", x"E8",
	x"E7", x"EE", x"F9", x"F7", x"F3", x"FA", x"02", x"06", x"03", x"FF", x"FB", x"FA",
	x"04", x"09", x"06", x"05", x"0A", x"11", x"10", x"0F", x"15", x"1A", x"14", x"0A",
	x"0C", x"16", x"17", x"0D", x"04", x"03", x"08", x"0A", x"08", x"0A", x"13", x"19",
	x"18", x"12", x"11", x"12", x"0E", x"0F", x"16", x"16", x"0F", x"09", x"08", x"0A",
	x"09", x"06", x"08", x"0D", x"0C", x"09", x"09", x"0D", x"0F", x"0A", x"03", x"FD",
	x"F6", x"F2", x"F8", x"FB", x"FE", x"02", x"FD", x"EE", x"E2", x"E5", x"F2", x"FA",
	x"F6", x"F0", x"F1", x"F4", x"ED", x"E7", x"F1", x"F9", x"F2", x"EF", x"F4", x"FC",
	x"02", x"05", x"07", x"09", x"06", x"FE", x"F4", x"F2", x"FA", x"09", x"13", x"0E",
	x"05", x"06", x"08", x"01", x"FC", x"03", x"0B", x"0D", x"0D", x"0C", x"04", x"F6",
	x"F1", x"F6", x"F6", x"F2", x"F8", x"00", x"FB", x"F2", x"F5", x"FE", x"03", x"FE",
	x"F6", x"EE", x"E9", x"E8", x"E8", x"EF", x"FC", x"FD", x"FA", x"FD", x"FE", x"F8",
	x"F2", x"F2", x"F7", x"F7", x"F4", x"F1", x"F2", x"F6", x"F4", x"F2", x"F3", x"EE",
	x"EA", x"EC", x"F2", x"F7", x"FA", x"F9", x"F3", x"EB", x"E9", x"ED", x"ED", x"E3",
	x"DF", x"E5", x"F1", x"FB", x"FB", x"FA", x"FB", x"F9", x"F8", x"00", x"09", x"0A",
	x"05", x"01", x"FF", x"FC", x"FA", x"FC", x"FE", x"FD", x"FC", x"FD", x"01", x"03",
	x"04", x"04", x"06", x"08", x"09", x"05", x"FF", x"FD", x"FF", x"01", x"FF", x"FC",
	x"FE", x"06", x"08", x"FB", x"F5", x"FD", x"01", x"FC", x"F9", x"00", x"0B", x"0C",
	x"0B", x"13", x"18", x"14", x"11", x"0F", x"0E", x"0C", x"07", x"09", x"13", x"19",
	x"13", x"0A", x"07", x"0E", x"1A", x"1C", x"1A", x"18", x"16", x"14", x"12", x"14",
	x"1A", x"18", x"0D", x"04", x"02", x"00", x"FF", x"01", x"02", x"03", x"08", x"0F",
	x"0D", x"06", x"0B", x"10", x"0F", x"0D", x"0E", x"0C", x"09", x"08", x"09", x"09",
	x"07", x"07", x"0B", x"0B", x"05", x"FE", x"FD", x"FA", x"ED", x"E6", x"ED", x"F4",
	x"F2", x"F0", x"F3", x"F5", x"F3", x"F0", x"F4", x"FA", x"FC", x"FB", x"F9", x"F9",
	x"FE", x"01", x"F9", x"EF", x"F1", x"FC", x"FD", x"F4", x"EF", x"F4", x"FB", x"F8",
	x"F0", x"EA", x"E6", x"E7", x"E6", x"E5", x"E7", x"EC", x"F1", x"F1", x"F0", x"F2",
	x"F3", x"F1", x"EE", x"ED", x"EF", x"F0", x"F0", x"F5", x"FA", x"F6", x"EB", x"E6",
	x"EC", x"F9", x"01", x"03", x"02", x"04", x"08", x"06", x"FE", x"F8", x"F2", x"F3",
	x"FF", x"05", x"01", x"02", x"08", x"0C", x"10", x"15", x"0D", x"04", x"05", x"04",
	x"05", x"0D", x"11", x"0E", x"09", x"02", x"FD", x"FF", x"03", x"07", x"0C", x"0C",
	x"06", x"FF", x"F7", x"F1", x"F2", x"F8", x"FE", x"01", x"FE", x"F8", x"FD", x"03",
	x"FC", x"F2", x"EC", x"E9", x"ED", x"F5", x"F6", x"EF", x"E9", x"E8", x"EB", x"EE",
	x"EB", x"E8", x"E8", x"EB", x"F0", x"F4", x"FD", x"0C", x"12", x"0E", x"07", x"02",
	x"00", x"05", x"0B", x"12", x"18", x"1C", x"19", x"11", x"10", x"13", x"15", x"16",
	x"15", x"12", x"0D", x"0E", x"12", x"0F", x"0F", x"1B", x"1E", x"13", x"0A", x"0D",
	x"11", x"0D", x"04", x"02", x"0A", x"13", x"12", x"0B", x"06", x"04", x"04", x"03",
	x"FF", x"FC", x"FB", x"01", x"06", x"00", x"FE", x"03", x"06", x"08", x"04", x"FE",
	x"FD", x"FD", x"FC", x"FC", x"00", x"03", x"FF", x"FC", x"01", x"05", x"05", x"09",
	x"0A", x"03", x"FE", x"02", x"04", x"00", x"00", x"01", x"FF", x"FB", x"FA", x"F9",
	x"F7", x"F6", x"F8", x"F6", x"EE", x"EE", x"F6", x"FA", x"F7", x"F3", x"F5", x"FB",
	x"01", x"03", x"02", x"02", x"05", x"05", x"04", x"02", x"03", x"06", x"04", x"FB",
	x"F9", x"03", x"0A", x"06", x"FA", x"F3", x"F2", x"F3", x"F4", x"F5", x"F8", x"FD",
	x"01", x"FE", x"F5", x"F2", x"F5", x"F8", x"FA", x"F8", x"F2", x"F2", x"FD", x"05",
	x"02", x"00", x"06", x"08", x"03", x"FF", x"02", x"08", x"0A", x"0A", x"0A", x"08",
	x"09", x"08", x"09", x"10", x"12", x"0C", x"03", x"F9", x"F4", x"F6", x"FA", x"FE",
	x"01", x"05", x"06", x"06", x"02", x"FE", x"FF", x"00", x"FE", x"00", x"02", x"FF",
	x"F8", x"F2", x"F2", x"F4", x"F6", x"F8", x"FF", x"05", x"01", x"F8", x"FA", x"02",
	x"08", x"08", x"06", x"08", x"0D", x"0D", x"0A", x"0A", x"0A", x"03", x"FE", x"FA",
	x"F8", x"FB", x"FC", x"F4", x"F0", x"F7", x"FC", x"F6", x"F1", x"F7", x"FC", x"F9",
	x"F4", x"F1", x"EF", x"ED", x"F0", x"F5", x"FB", x"02", x"03", x"FE", x"F7", x"F5",
	x"F5", x"F4", x"F1", x"E9", x"E6", x"E9", x"ED", x"F0", x"F0", x"F3", x"F8", x"FD",
	x"FD", x"F4", x"EA", x"E9", x"F2", x"FC", x"FE", x"FD", x"01", x"02", x"00", x"01",
	x"00", x"FE", x"02", x"09", x"0E", x"09", x"02", x"05", x"0D", x"12", x"11", x"0F",
	x"0C", x"0D", x"14", x"17", x"13", x"0E", x"09", x"08", x"0F", x"18", x"1E", x"1C",
	x"19", x"16", x"15", x"16", x"12", x"08", x"08", x"10", x"12", x"0B", x"06", x"05",
	x"03", x"FA", x"F2", x"EF", x"F0", x"F2", x"F1", x"F2", x"F6", x"F8", x"F3", x"ED",
	x"EF", x"F7", x"FF", x"FF", x"FC", x"FE", x"FF", x"FB", x"F9", x"01", x"07", x"05",
	x"00", x"FF", x"04", x"07", x"06", x"06", x"0A", x"0F", x"0E", x"0D", x"0F", x"12",
	x"15", x"14", x"0E", x"07", x"06", x"09", x"08", x"04", x"06", x"0B", x"10", x"0F",
	x"06", x"01", x"04", x"06", x"01", x"FA", x"FF", x"0A", x"07", x"F9", x"F4", x"FC",
	x"05", x"04", x"FA", x"F3", x"EE", x"ED", x"EF", x"F5", x"F8", x"FB", x"FF", x"FE",
	x"FC", x"FA", x"F7", x"F6", x"F9", x"FC", x"FD", x"FD", x"FB", x"F8", x"F8", x"F6",
	x"F7", x"F9", x"F9", x"F3", x"EE", x"F0", x"F6", x"F9", x"F6", x"F2", x"F1", x"F1",
	x"F2", x"F3", x"EF", x"EC", x"EE", x"F3", x"F6", x"F8", x"F9", x"F8", x"F4", x"F2",
	x"F8", x"02", x"08", x"07", x"FE", x"F2", x"EF", x"F6", x"FB", x"FC", x"FD", x"FD",
	x"FA", x"F0", x"E8", x"EA", x"F0", x"F2", x"F2", x"F4", x"F3", x"EF", x"F1", x"F6",
	x"FA", x"FD", x"F9", x"F2", x"F5", x"FC", x"FF", x"05", x"11", x"19", x"11", x"03",
	x"05", x"0E", x"0B", x"07", x"08", x"09", x"0B", x"07", x"05", x"0A", x"08", x"05",
	x"0A", x"0F", x"12", x"10", x"0A", x"0A", x"11", x"18", x"19", x"16", x"16", x"13",
	x"0D", x"0B", x"10", x"12", x"09", x"03", x"03", x"00", x"F9", x"F7", x"FD", x"04",
	x"0A", x"07", x"FD", x"F6", x"F9", x"02", x"0B", x"0B", x"04", x"01", x"01", x"00",
	x"04", x"09", x"0D", x"08", x"01", x"03", x"09", x"0E", x"0D", x"0D", x"14", x"1C",
	x"1A", x"15", x"12", x"14", x"15", x"0D", x"03", x"02", x"04", x"06", x"05", x"02",
	x"00", x"FC", x"FA", x"FA", x"F8", x"F4", x"F0", x"F0", x"F2", x"F9", x"00", x"FE",
	x"F5", x"F0", x"F2", x"F7", x"FC", x"01", x"01", x"FB", x"F7", x"F7", x"F4", x"EC",
	x"EB", x"EE", x"EF", x"EE", x"F2", x"F8", x"FC", x"FA", x"F8", x"F7", x"EE", x"E3",
	x"E0", x"E6", x"EF", x"F2", x"F6", x"FB", x"FE", x"00", x"00", x"00", x"04", x"0C",
	x"10", x"0D", x"0A", x"0C", x"11", x"10", x"09", x"04", x"FF", x"FC", x"FE", x"FF",
	x"FB", x"F9", x"FF", x"06", x"04", x"03", x"07", x"0A", x"0B", x"06", x"FE", x"FB",
	x"FE", x"FE", x"F8", x"F9", x"FF", x"FF", x"F9", x"F5", x"F5", x"F6", x"F4", x"F2",
	x"F1", x"F3", x"F2", x"EE", x"EC", x"EC", x"F1", x"F4", x"F3", x"F6", x"FD", x"01",
	x"FF", x"FA", x"F7", x"F8", x"FB", x"FF", x"01", x"01", x"03", x"04", x"00", x"FF",
	x"03", x"07", x"01", x"F9", x"F9", x"00", x"06", x"08", x"0A", x"0D", x"0B", x"08",
	x"0C", x"11", x"12", x"11", x"10", x"10", x"0F", x"0E", x"0F", x"0E", x"06", x"02",
	x"FE", x"F5", x"F2", x"F6", x"F7", x"F4", x"F7", x"FD", x"02", x"06", x"09", x"09",
	x"0A", x"0C", x"0E", x"0F", x"09", x"02", x"03", x"04", x"01", x"FE", x"02", x"06",
	x"03", x"FF", x"FC", x"F7", x"F4", x"FB", x"01", x"00", x"FA", x"F4", x"F5", x"FC",
	x"03", x"05", x"06", x"0E", x"12", x"0A", x"FE", x"FB", x"FD", x"FB", x"F9", x"F8",
	x"F7", x"F8", x"F9", x"F4", x"F2", x"F6", x"FA", x"F8", x"F7", x"F9", x"FB", x"F9",
	x"F5", x"F7", x"FD", x"02", x"04", x"06", x"03", x"FB", x"F4", x"F5", x"FA", x"FB",
	x"FA", x"F9", x"F8", x"F9", x"FD", x"00", x"02", x"FF", x"F9", x"FA", x"01", x"05",
	x"05", x"05", x"03", x"FF", x"FD", x"F8", x"F6", x"FC", x"FE", x"F6", x"F0", x"F7",
	x"05", x"0D", x"0A", x"04", x"04", x"06", x"05", x"06", x"07", x"07", x"09", x"08",
	x"04", x"00", x"03", x"07", x"09", x"08", x"09", x"0D", x"0D", x"0B", x"07", x"08",
	x"0A", x"09", x"08", x"09", x"08", x"04", x"04", x"04", x"04", x"06", x"03", x"FC",
	x"F4", x"F2", x"F5", x"F8", x"FA", x"FB", x"F9", x"F9", x"00", x"05", x"04", x"02",
	x"04", x"07", x"08", x"07", x"04", x"03", x"03", x"02", x"02", x"02", x"03", x"03",
	x"01", x"01", x"00", x"FC", x"FB", x"FF", x"FD", x"F7", x"F9", x"FB", x"FA", x"F7",
	x"F9", x"FE", x"03", x"02", x"FA", x"F7", x"FB", x"FD", x"F7", x"ED", x"EE", x"F5",
	x"FA", x"F6", x"F4", x"F4", x"F1", x"ED", x"EC", x"EA", x"EA", x"ED", x"EF", x"F1",
	x"F2", x"F1", x"EB", x"EB", x"F5", x"FB", x"FB", x"01", x"08", x"08", x"FD", x"F4",
	x"F6", x"FA", x"F9", x"FE", x"07", x"0A", x"04", x"FF", x"03", x"09", x"08", x"06",
	x"06", x"06", x"04", x"05", x"0B", x"0D", x"09", x"09", x"08", x"03", x"00", x"00",
	x"02", x"03", x"02", x"01", x"00", x"00", x"02", x"04", x"02", x"00", x"FF", x"04",
	x"0A", x"09", x"08", x"08", x"09", x"08", x"08", x"09", x"07", x"03", x"FA", x"F5",
	x"F8", x"FC", x"FE", x"FC", x"F7", x"F5", x"F6", x"FC", x"01", x"FF", x"FD", x"FF",
	x"FF", x"FD", x"FA", x"FD", x"00", x"00", x"03", x"08", x"0C", x"09", x"03", x"FE",
	x"FC", x"FD", x"00", x"07", x"0C", x"0D", x"0B", x"0D", x"0F", x"0C", x"08", x"08",
	x"09", x"09", x"05", x"04", x"03", x"00", x"FE", x"FD", x"FD", x"FF", x"05", x"0C",
	x"0A", x"05", x"03", x"06", x"05", x"FC", x"F8", x"FC", x"FF", x"F6", x"F2", x"FC",
	x"05", x"06", x"01", x"FC", x"FE", x"02", x"02", x"03", x"07", x"03", x"FB", x"FA",
	x"01", x"07", x"06", x"03", x"03", x"FF", x"F7", x"F8", x"FF", x"04", x"05", x"04",
	x"00", x"FC", x"F9", x"F9", x"FA", x"FD", x"FC", x"F4", x"EC", x"EE", x"F6", x"F9",
	x"F6", x"F0", x"ED", x"ED", x"EE", x"F0", x"F5", x"FC", x"02", x"02", x"FC", x"F6",
	x"F4", x"F5", x"F5", x"F4", x"F3", x"F3", x"F5", x"FA", x"FC", x"FC", x"FF", x"00",
	x"FE", x"FB", x"FF", x"06", x"07", x"03", x"FE", x"FC", x"FD", x"FD", x"FB", x"FB",
	x"01", x"06", x"04", x"FF", x"FF", x"03", x"06", x"04", x"00", x"00", x"04", x"05",
	x"02", x"04", x"06", x"02", x"F9", x"F7", x"FD", x"05", x"07", x"03", x"00", x"02",
	x"05", x"02", x"FF", x"FE", x"00", x"01", x"FF", x"00", x"05", x"04", x"00", x"FD",
	x"01", x"04", x"01", x"FD", x"FF", x"04", x"07", x"08", x"06", x"03", x"07", x"0D",
	x"11", x"0E", x"0C", x"0C", x"09", x"08", x"0B", x"08", x"01", x"00", x"04", x"07",
	x"07", x"04", x"00", x"00", x"01", x"02", x"06", x"09", x"06", x"01", x"FE", x"FF",
	x"04", x"05", x"03", x"04", x"07", x"05", x"01", x"FB", x"F8", x"FF", x"04", x"FD",
	x"F3", x"F1", x"F8", x"00", x"FC", x"F2", x"EE", x"F1", x"F4", x"F2", x"F1", x"F1",
	x"F0", x"ED", x"EB", x"F0", x"FC", x"00", x"FD", x"FA", x"FC", x"01", x"03", x"03",
	x"05", x"07", x"04", x"FF", x"FE", x"01", x"03", x"03", x"01", x"00", x"03", x"06",
	x"08", x"09", x"06", x"01", x"F8", x"F0", x"F1", x"F9", x"F8", x"F3", x"F7", x"02",
	x"06", x"01", x"01", x"06", x"05", x"00", x"FB", x"FB", x"FC", x"F9", x"F7", x"FD",
	x"01", x"FE", x"F9", x"F6", x"F4", x"F5", x"F9", x"FD", x"FD", x"FC", x"FB", x"FA",
	x"FB", x"FD", x"FD", x"FD", x"00", x"FF", x"FD", x"00", x"04", x"05", x"02", x"FD",
	x"FD", x"FF", x"FD", x"FB", x"FB", x"00", x"04", x"03", x"FF", x"FD", x"FE", x"03",
	x"07", x"06", x"02", x"01", x"00", x"03", x"04", x"00", x"01", x"06", x"0A", x"0A",
	x"08", x"04", x"FF", x"FF", x"03", x"04", x"FF", x"FB", x"FD", x"01", x"01", x"FF",
	x"FF", x"04", x"08", x"06", x"FF", x"FB", x"FC", x"FE", x"FF", x"FF", x"02", x"06",
	x"08", x"07", x"04", x"04", x"05", x"02", x"FF", x"FF", x"01", x"00", x"00", x"FE",
	x"FC", x"01", x"09", x"0B", x"06", x"FE", x"FE", x"06", x"0B", x"0C", x"0A", x"08",
	x"05", x"01", x"FE", x"00", x"04", x"05", x"03", x"FF", x"FB", x"FB", x"01", x"08",
	x"09", x"01", x"FB", x"F8", x"F7", x"F7", x"F8", x"F8", x"F9", x"F9", x"F8", x"F6",
	x"F5", x"F4", x"F6", x"F7", x"F7", x"F8", x"F6", x"F2", x"EF", x"ED", x"EE", x"EF",
	x"EF", x"EF", x"EF", x"EF", x"EE", x"ED", x"EF", x"F5", x"F7", x"F8", x"F8", x"F7",
	x"F9", x"FA", x"FC", x"00", x"05", x"07", x"06", x"06", x"04", x"01", x"01", x"02",
	x"06", x"08", x"07", x"06", x"07", x"09", x"05", x"05", x"0A", x"0D", x"0B", x"09",
	x"06", x"03", x"05", x"0C", x"0B", x"05", x"00", x"FC", x"FD", x"FF", x"02", x"01",
	x"00", x"00", x"FE", x"FC", x"FD", x"00", x"01", x"05", x"0C", x"0E", x"09", x"08",
	x"0C", x"0D", x"0A", x"0A", x"0B", x"07", x"00", x"00", x"0A", x"11", x"0E", x"07",
	x"02", x"01", x"03", x"06", x"07", x"07", x"07", x"07", x"07", x"0B", x"0D", x"0A",
	x"08", x"08", x"07", x"04", x"02", x"03", x"08", x"0B", x"09", x"03", x"FD", x"FD",
	x"04", x"0A", x"0A", x"06", x"00", x"FC", x"FC", x"FC", x"FC", x"FE", x"FB", x"F5",
	x"EF", x"EE", x"F1", x"F4", x"F3", x"F0", x"F2", x"F3", x"F1", x"F2", x"F4", x"F5",
	x"F5", x"F4", x"F5", x"F6", x"F6", x"F7", x"F7", x"F7", x"F8", x"FA", x"FC", x"F8",
	x"F3", x"F4", x"F9", x"FC", x"F9", x"F8", x"FB", x"FF", x"01", x"02", x"02", x"04",
	x"05", x"07", x"06", x"06", x"04", x"01", x"02", x"02", x"FF", x"FF", x"00", x"03",
	x"00", x"FC", x"FD", x"FC", x"F9", x"F8", x"F9", x"F6", x"F6", x"F7", x"F7", x"F9",
	x"FA", x"FB", x"FC", x"FA", x"F9", x"FA", x"FC", x"FD", x"FE", x"FE", x"FC", x"FC",
	x"FE", x"FF", x"FC", x"FA", x"FA", x"FC", x"FE", x"FD", x"FA", x"F8", x"FA", x"FE",
	x"FD", x"FC", x"FD", x"FF", x"00", x"01", x"05", x"09", x"0A", x"09", x"09", x"09",
	x"08", x"06", x"07", x"0C", x"0D", x"0B", x"09", x"0A", x"0B", x"0C", x"0C", x"09",
	x"07", x"07", x"04", x"02", x"03", x"06", x"07", x"07", x"05", x"01", x"FF", x"04",
	x"08", x"06", x"01", x"FC", x"FD", x"02", x"03", x"FF", x"FE", x"00", x"00", x"FE",
	x"FB", x"F9", x"FA", x"F9", x"F7", x"F6", x"F6", x"F4", x"F5", x"F7", x"F8", x"FB",
	x"04", x"0A", x"0B", x"09", x"08", x"08", x"07", x"05", x"04", x"05", x"05", x"06",
	x"04", x"04", x"06", x"09", x"0D", x"0F", x"0D", x"0A", x"06", x"03", x"04", x"06",
	x"05", x"03", x"02", x"01", x"FD", x"FB", x"FC", x"FF", x"FF", x"FF", x"FF", x"FC",
	x"F9", x"F7", x"F4", x"F4", x"F7", x"F9", x"F5", x"F2", x"F3", x"F4", x"F2", x"F1",
	x"F3", x"F5", x"F4", x"F0", x"EE", x"F1", x"F5", x"F5", x"F4", x"F6", x"F8", x"F8",
	x"F5", x"F5", x"FB", x"FD", x"FA", x"F8", x"FA", x"FD", x"FB", x"FC", x"03", x"07",
	x"05", x"03", x"04", x"04", x"06", x"08", x"07", x"07", x"06", x"04", x"02", x"FF",
	x"FD", x"FB", x"F9", x"F9", x"FD", x"01", x"03", x"01", x"FE", x"FF", x"02", x"03",
	x"05", x"05", x"03", x"03", x"05", x"02", x"FE", x"FF", x"02", x"03", x"01", x"FF",
	x"FD", x"FB", x"FE", x"03", x"03", x"01", x"00", x"01", x"FE", x"FC", x"FE", x"00",
	x"03", x"07", x"08", x"07", x"05", x"05", x"03", x"03", x"04", x"06", x"05", x"03",
	x"04", x"07", x"0C", x"0F", x"0D", x"0B", x"0E", x"10", x"0C", x"06", x"05", x"07",
	x"06", x"05", x"04", x"02", x"FE", x"FA", x"F9", x"FC", x"FF", x"FC", x"F7", x"F6",
	x"F7", x"F7", x"F8", x"FD", x"01", x"FD", x"F5", x"F4", x"FC", x"03", x"02", x"FD",
	x"F9", x"F7", x"F7", x"F8", x"F6", x"F7", x"FB", x"FC", x"FA", x"F7", x"F4", x"F3",
	x"F3", x"F9", x"02", x"04", x"FF", x"FE", x"01", x"03", x"02", x"02", x"06", x"08",
	x"04", x"00", x"01", x"07", x"08", x"02", x"00", x"03", x"01", x"FC", x"FA", x"FC",
	x"00", x"FE", x"FB", x"FE", x"02", x"00", x"FB", x"FB", x"FC", x"FC", x"FD", x"FB",
	x"FB", x"FD", x"FD", x"F7", x"F4", x"FA", x"01", x"02", x"00", x"00", x"01", x"FE",
	x"FB", x"FD", x"00", x"FD", x"F8", x"F7", x"FA", x"FD", x"FC", x"FB", x"FC", x"FE",
	x"FE", x"FC", x"F9", x"F8", x"F9", x"FC", x"FD", x"FE", x"FF", x"03", x"05", x"04",
	x"02", x"05", x"08", x"08", x"05", x"05", x"09", x"0A", x"08", x"06", x"09", x"0D",
	x"0C", x"08", x"04", x"01", x"01", x"05", x"08", x"06", x"06", x"0A", x"0B", x"09",
	x"09", x"0B", x"09", x"08", x"0B", x"0A", x"04", x"01", x"02", x"03", x"01", x"FE",
	x"FD", x"FE", x"FE", x"F9", x"F4", x"F4", x"F7", x"FB", x"F9", x"F7", x"FC", x"02",
	x"00", x"FE", x"02", x"08", x"0A", x"06", x"01", x"02", x"03", x"02", x"01", x"03",
	x"05", x"04", x"FF", x"FB", x"F9", x"F9", x"FA", x"FD", x"FD", x"FA", x"F8", x"FC",
	x"00", x"FE", x"FB", x"FC", x"FF", x"FF", x"02", x"03", x"FF", x"FB", x"F8", x"F9",
	x"FA", x"F9", x"F7", x"F6", x"F6", x"F7", x"F8", x"F9", x"FA", x"FC", x"FE", x"FF",
	x"FE", x"FA", x"FA", x"FB", x"FA", x"FA", x"FB", x"FD", x"FB", x"F9", x"FA", x"FC",
	x"FB", x"F7", x"F5", x"F8", x"FF", x"01", x"FD", x"FC", x"01", x"03", x"02", x"00",
	x"FE", x"FE", x"01", x"04", x"03", x"01", x"00", x"FE", x"FC", x"FB", x"FD", x"FC",
	x"F9", x"FA", x"FC", x"FD", x"FE", x"FD", x"FD", x"02", x"05", x"02", x"FF", x"01",
	x"05", x"09", x"0A", x"0C", x"0E", x"0E", x"0F", x"10", x"0D", x"09", x"0B", x"0C",
	x"08", x"02", x"FF", x"FE", x"00", x"00", x"FE", x"FF", x"FF", x"FF", x"FF", x"03",
	x"08", x"05", x"01", x"01", x"03", x"05", x"05", x"03", x"00", x"01", x"05", x"07",
	x"06", x"05", x"07", x"07", x"01", x"FC", x"FB", x"F8", x"F5", x"F7", x"FA", x"FC",
	x"FD", x"FE", x"FF", x"01", x"02", x"00", x"00", x"01", x"02", x"FF", x"F9", x"F9",
	x"FF", x"05", x"05", x"02", x"03", x"04", x"01", x"FD", x"FB", x"FB", x"FB", x"FC",
	x"FB", x"F9", x"FC", x"00", x"03", x"02", x"FF", x"FF", x"01", x"03", x"00", x"FE",
	x"FB", x"F9", x"F9", x"F9", x"F7", x"F6", x"F8", x"F8", x"F8", x"FB", x"FB", x"F8",
	x"F7", x"FA", x"00", x"01", x"FD", x"FC", x"00", x"03", x"01", x"FF", x"02", x"00",
	x"FB", x"F9", x"FA", x"FA", x"F9", x"F7", x"F7", x"FB", x"FA", x"F4", x"F4", x"F9",
	x"FB", x"FA", x"FB", x"02", x"06", x"00", x"FB", x"FE", x"01", x"FF", x"FB", x"FD",
	x"02", x"03", x"04", x"07", x"0A", x"06", x"00", x"FD", x"FA", x"F8", x"F8", x"F8",
	x"F9", x"FE", x"01", x"FE", x"FB", x"FA", x"F9", x"F9", x"FD", x"01", x"00", x"FE",
	x"FF", x"01", x"03", x"05", x"07", x"06", x"03", x"01", x"01", x"02", x"04", x"06",
	x"06", x"05", x"03", x"03", x"05", x"08", x"07", x"06", x"06", x"08", x"09", x"07",
	x"03", x"02", x"05", x"06", x"04", x"03", x"03", x"03", x"03", x"00", x"FE", x"02",
	x"07", x"0A", x"0C", x"0D", x"0A", x"02", x"00", x"03", x"07", x"09", x"06", x"05",
	x"04", x"03", x"03", x"04", x"04", x"04", x"01", x"FD", x"FA", x"FB", x"FE", x"03",
	x"05", x"03", x"FC", x"F8", x"FB", x"FF", x"02", x"01", x"FE", x"FB", x"F5", x"F3",
	x"F5", x"F6", x"F7", x"F8", x"FA", x"FC", x"F9", x"F7", x"F9", x"FC", x"FC", x"F8",
	x"F6", x"F6", x"F7", x"FA", x"FD", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE", x"FE",
	x"FA", x"F7", x"F8", x"FA", x"FB", x"FD", x"FE", x"FF", x"FF", x"00", x"02", x"01",
	x"00", x"02", x"01", x"FD", x"FB", x"FB", x"FD", x"FF", x"00", x"00", x"02", x"03",
	x"03", x"FE", x"F9", x"FA", x"FC", x"FE", x"FE", x"FD", x"FD", x"00", x"FA", x"F2",
	x"F1", x"F7", x"F9", x"F7", x"F5", x"F5", x"F9", x"FF", x"03", x"02", x"FF", x"00",
	x"02", x"02", x"FF", x"FE", x"02", x"04", x"03", x"01", x"02", x"05", x"05", x"06",
	x"08", x"0B", x"0E", x"0C", x"07", x"05", x"08", x"0C", x"0D", x"0B", x"09", x"0C",
	x"0C", x"0B", x"0A", x"0A", x"09", x"04", x"00", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FF", x"01", x"00", x"FE", x"FD", x"01", x"05", x"04", x"01", x"00", x"01",
	x"00", x"FF", x"02", x"03", x"00", x"FB", x"FA", x"FE", x"FF", x"FC", x"F9", x"F8",
	x"FC", x"00", x"00", x"FD", x"FD", x"FF", x"FF", x"FA", x"F4", x"F5", x"FD", x"04",
	x"04", x"01", x"FF", x"FE", x"FF", x"00", x"FE", x"FF", x"00", x"02", x"01", x"01",
	x"01", x"02", x"02", x"FF", x"FE", x"00", x"01", x"00", x"FE", x"FE", x"00", x"04",
	x"06", x"04", x"02", x"03", x"06", x"06", x"00", x"F8", x"F3", x"F4", x"F8", x"F9",
	x"F7", x"F7", x"F8", x"F8", x"F6", x"F4", x"F2", x"F4", x"F6", x"F8", x"FA", x"F8",
	x"F8", x"FC", x"00", x"02", x"04", x"03", x"FF", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"FF", x"FC", x"FB", x"FC", x"FC",
	x"FD", x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FA", x"F9", x"FD", x"01", x"02",
	x"01", x"FF", x"00", x"02", x"03", x"02", x"FF", x"FE", x"FE", x"FB", x"F9", x"FB",
	x"FF", x"04", x"09", x"08", x"03", x"FE", x"FF", x"04", x"06", x"03", x"03", x"08",
	x"0A", x"06", x"02", x"03", x"06", x"05", x"01", x"03", x"09", x"08", x"04", x"01",
	x"01", x"04", x"05", x"03", x"00", x"FD", x"FE", x"02", x"07", x"08", x"09", x"09",
	x"05", x"01", x"04", x"07", x"05", x"02", x"01", x"03", x"02", x"FF", x"FF", x"00",
	x"02", x"02", x"FE", x"FB", x"FA", x"F8", x"F8", x"F9", x"FB", x"FA", x"F9", x"F8",
	x"F5", x"F5", x"F7", x"F7", x"F4", x"F3", x"F3", x"F3", x"F2", x"F3", x"F6", x"F7",
	x"F6", x"F8", x"FC", x"FB", x"F6", x"F6", x"FD", x"01", x"FD", x"F8", x"F7", x"F8",
	x"FB", x"FE", x"FF", x"00", x"00", x"02", x"06", x"06", x"05", x"05", x"05", x"02",
	x"00", x"FF", x"00", x"02", x"04", x"06", x"06", x"02", x"00", x"01", x"01", x"FF",
	x"FE", x"FC", x"FB", x"FC", x"FD", x"FE", x"FE", x"FD", x"FD", x"FE", x"FC", x"FB",
	x"FB", x"FD", x"FD", x"FB", x"FB", x"FD", x"02", x"02", x"FA", x"F4", x"F6", x"FA",
	x"FC", x"FC", x"00", x"06", x"07", x"04", x"00", x"00", x"02", x"05", x"05", x"05",
	x"06", x"0A", x"0D", x"0C", x"0C", x"12", x"14", x"0E", x"09", x"0A", x"0F", x"0F",
	x"0B", x"08", x"08", x"0A", x"08", x"04", x"06", x"0A", x"0A", x"07", x"05", x"04",
	x"01", x"FE", x"FD", x"FD", x"FD", x"FD", x"00", x"02", x"01", x"FF", x"FD", x"FD",
	x"FD", x"FC", x"F9", x"F6", x"F5", x"F5", x"F6", x"F7", x"F8", x"FC", x"FF", x"FE",
	x"FB", x"FC", x"FE", x"FD", x"FB", x"FA", x"FD", x"01", x"FF", x"FC", x"FD", x"FF",
	x"FD", x"F9", x"F8", x"FA", x"FC", x"FE", x"00", x"00", x"00", x"FF", x"FF", x"01",
	x"03", x"05", x"06", x"07", x"0A", x"08", x"03", x"00", x"01", x"02", x"00", x"FE",
	x"FE", x"FD", x"FE", x"01", x"00", x"FC", x"F9", x"F7", x"F6", x"F5", x"F2", x"F2",
	x"F6", x"F8", x"F5", x"F5", x"F7", x"F8", x"F8", x"F7", x"F6", x"F6", x"F8", x"FA",
	x"F9", x"F7", x"F9", x"FB", x"FC", x"FC", x"FC", x"FF", x"02", x"02", x"FF", x"FB",
	x"FA", x"FB", x"FB", x"FA", x"F8", x"F7", x"F7", x"F9", x"FC", x"00", x"03", x"04",
	x"03", x"00", x"FD", x"FD", x"FF", x"FF", x"FE", x"FD", x"FB", x"FA", x"00", x"04",
	x"04", x"05", x"07", x"07", x"02", x"FF", x"01", x"06", x"05", x"00", x"FE", x"01",
	x"03", x"04", x"02", x"00", x"04", x"08", x"08", x"05", x"06", x"0A", x"0B", x"08",
	x"03", x"FD", x"FE", x"00", x"02", x"05", x"09", x"06", x"01", x"FF", x"01", x"04",
	x"06", x"08", x"09", x"09", x"07", x"04", x"03", x"07", x"0A", x"0B", x"0B", x"0B",
	x"0A", x"0A", x"0B", x"0C", x"0C", x"0A", x"09", x"09", x"08", x"08", x"08", x"07",
	x"05", x"FF", x"F8", x"F5", x"F5", x"FA", x"FE", x"FE", x"FC", x"FB", x"FB", x"F9",
	x"F7", x"F7", x"F7", x"F8", x"F8", x"FA", x"FA", x"F9", x"F9", x"F9", x"F7", x"F8",
	x"FC", x"FC", x"FB", x"FD", x"00", x"02", x"00", x"FD", x"FB", x"FD", x"FE", x"FE",
	x"FC", x"F8", x"F6", x"F7", x"FA", x"FA", x"FA", x"FB", x"FA", x"FA", x"FC", x"FF",
	x"03", x"06", x"06", x"03", x"01", x"00", x"FD", x"FD", x"FF", x"01", x"FE", x"FB",
	x"FA", x"FC", x"FC", x"FB", x"FA", x"F8", x"F6", x"F4", x"F3", x"F5", x"FA", x"FD",
	x"FC", x"FA", x"FB", x"FB", x"F9", x"F8", x"FB", x"01", x"02", x"00", x"FD", x"FD",
	x"FF", x"FD", x"FC", x"01", x"09", x"0A", x"05", x"00", x"FF", x"00", x"02", x"02",
	x"00", x"02", x"04", x"00", x"FA", x"FE", x"08", x"0A", x"07", x"06", x"09", x"09",
	x"05", x"03", x"06", x"09", x"07", x"05", x"03", x"04", x"05", x"02", x"00", x"FE",
	x"FB", x"FA", x"FB", x"FF", x"02", x"00", x"FF", x"02", x"04", x"02", x"01", x"03",
	x"04", x"00", x"FB", x"FC", x"01", x"01", x"FB", x"FA", x"FD", x"01", x"00", x"FD",
	x"FD", x"FD", x"FB", x"F8", x"F5", x"F7", x"FC", x"FF", x"FE", x"00", x"04", x"02",
	x"FC", x"F9", x"FB", x"FC", x"FD", x"FD", x"FD", x"FD", x"FE", x"02", x"03", x"00",
	x"00", x"01", x"00", x"00", x"FE", x"FD", x"00", x"04", x"05", x"03", x"05", x"05",
	x"04", x"03", x"00", x"FE", x"FF", x"02", x"02", x"FE", x"FD", x"FF", x"FF", x"F9",
	x"F6", x"F9", x"FF", x"01", x"FF", x"FE", x"FF", x"FF", x"FB", x"F6", x"F4", x"F5",
	x"F6", x"FA", x"FF", x"01", x"FF", x"01", x"06", x"05", x"00", x"FD", x"FF", x"FF",
	x"FB", x"F9", x"FA", x"FD", x"00", x"03", x"03", x"02", x"03", x"06", x"04", x"FE",
	x"FB", x"FA", x"FA", x"FC", x"01", x"05", x"06", x"03", x"01", x"00", x"01", x"00",
	x"FD", x"FE", x"02", x"06", x"08", x"07", x"02", x"FE", x"FD", x"FC", x"FC", x"00",
	x"01", x"01", x"03", x"05", x"05", x"06", x"07", x"06", x"04", x"05", x"06", x"05",
	x"06", x"0B", x"0D", x"09", x"05", x"06", x"09", x"07", x"04", x"06", x"08", x"04",
	x"01", x"01", x"05", x"07", x"04", x"02", x"02", x"02", x"05", x"08", x"05", x"02",
	x"02", x"06", x"06", x"04", x"03", x"03", x"00", x"FA", x"F7", x"F9", x"FC", x"FB",
	x"F9", x"F6", x"F5", x"F7", x"FB", x"FC", x"FB", x"F9", x"F7", x"F7", x"F6", x"F5",
	x"F4", x"F5", x"F5", x"F7", x"F9", x"F9", x"F7", x"F7", x"F8", x"F8", x"F4", x"F3",
	x"F6", x"FB", x"00", x"04", x"03", x"FB", x"F9", x"FC", x"FE", x"02", x"05", x"06",
	x"03", x"FD", x"FB", x"FC", x"FF", x"FE", x"FA", x"F8", x"FA", x"FD", x"FE", x"01",
	x"02", x"00", x"FE", x"FE", x"FD", x"FC", x"FA", x"F8", x"F7", x"F8", x"FC", x"00",
	x"01", x"FF", x"FD", x"FC", x"FA", x"F7", x"F6", x"F9", x"F8", x"F5", x"F5", x"F7",
	x"F9", x"F9", x"F8", x"F8", x"FA", x"FC", x"00", x"05", x"09", x"0B", x"09", x"07",
	x"06", x"05", x"02", x"FF", x"FF", x"00", x"04", x"09", x"0C", x"0A", x"06", x"05",
	x"05", x"03", x"FE", x"FE", x"03", x"05", x"02", x"FF", x"FF", x"03", x"06", x"06",
	x"07", x"09", x"08", x"03", x"FF", x"02", x"06", x"03", x"00", x"01", x"06", x"09",
	x"07", x"07", x"08", x"08", x"05", x"03", x"04", x"05", x"06", x"05", x"04", x"04",
	x"06", x"07", x"05", x"00", x"FC", x"FB", x"FF", x"03", x"05", x"09", x"0C", x"09",
	x"03", x"FE", x"FE", x"01", x"03", x"03", x"02", x"03", x"04", x"03", x"03", x"05",
	x"06", x"04", x"FF", x"FD", x"FD", x"FD", x"FE", x"01", x"02", x"01", x"00", x"FC",
	x"FB", x"FF", x"01", x"FD", x"FB", x"FC", x"F9", x"F4", x"F2", x"F4", x"F6", x"F7",
	x"FA", x"FC", x"FF", x"00", x"FC", x"F8", x"F8", x"F9", x"F8", x"FB", x"00", x"04",
	x"05", x"02", x"FC", x"F9", x"FC", x"FE", x"FF", x"00", x"FE", x"FA", x"F7", x"F7",
	x"FA", x"FD", x"FD", x"FB", x"FD", x"FF", x"FC", x"FB", x"FB", x"FC", x"FB", x"FB",
	x"FD", x"FD", x"FB", x"FA", x"FB", x"FC", x"FA", x"F6", x"F4", x"F4", x"F2", x"F0",
	x"F1", x"F5", x"F9", x"FA", x"FA", x"FC", x"FD", x"FD", x"FE", x"01", x"02", x"FD",
	x"F9", x"FB", x"FD", x"FF", x"00", x"02", x"01", x"00", x"02", x"04", x"00", x"FC",
	x"FD", x"FE", x"FC", x"FB", x"01", x"0B", x"10", x"0F", x"0F", x"10", x"11", x"10",
	x"0B", x"0A", x"0C", x"0F", x"0F", x"0E", x"0A", x"06", x"06", x"05", x"FF", x"FD",
	x"FF", x"FF", x"FC", x"FD", x"FF", x"FF", x"FE", x"FE", x"00", x"02", x"02", x"00",
	x"02", x"05", x"04", x"00", x"FE", x"FF", x"FF", x"FD", x"FC", x"FB", x"F9", x"F7",
	x"F8", x"FA", x"F9", x"F7", x"F7", x"F7", x"F6", x"F5", x"F5", x"F7", x"F8", x"F8",
	x"F9", x"FB", x"FC", x"FB", x"FC", x"FD", x"FE", x"FE", x"FF", x"00", x"04", x"06",
	x"04", x"01", x"02", x"03", x"01", x"FE", x"FF", x"03", x"03", x"FF", x"FE", x"01",
	x"04", x"05", x"03", x"05", x"06", x"04", x"03", x"04", x"03", x"00", x"FE", x"FF",
	x"00", x"03", x"03", x"02", x"03", x"00", x"FC", x"FC", x"FC", x"FA", x"F9", x"FA",
	x"FB", x"FA", x"F8", x"F8", x"FA", x"FC", x"FF", x"01", x"01", x"FB", x"F7", x"F7",
	x"FB", x"FC", x"FD", x"00", x"01", x"00", x"FE", x"FE", x"02", x"03", x"03", x"03",
	x"04", x"06", x"07", x"06", x"09", x"10", x"13", x"0F", x"08", x"07", x"08", x"07",
	x"04", x"05", x"04", x"01", x"00", x"FE", x"FD", x"FC", x"FD", x"00", x"02", x"01",
	x"FD", x"F9", x"F8", x"FB", x"FE", x"FE", x"FD", x"FD", x"FF", x"02", x"01", x"00",
	x"01", x"03", x"03", x"02", x"04", x"07", x"05", x"04", x"03", x"03", x"04", x"06",
	x"07", x"06", x"04", x"03", x"01", x"00", x"00", x"FE", x"FD", x"FD", x"FE", x"FF",
	x"00", x"03", x"06", x"04", x"01", x"FE", x"FF", x"02", x"05", x"02", x"FE", x"FE",
	x"01", x"01", x"00", x"01", x"03", x"01", x"FC", x"F9", x"FA", x"FA", x"F9", x"F9",
	x"FA", x"F9", x"F7", x"F3", x"F3", x"F6", x"F9", x"FC", x"FD", x"F9", x"F5", x"F2",
	x"F0", x"F2", x"F7", x"F9", x"FB", x"FB", x"F8", x"F5", x"F3", x"F3", x"FA", x"03",
	x"04", x"FF", x"FB", x"FA", x"FB", x"FB", x"FF", x"06", x"08", x"04", x"FF", x"FF",
	x"FF", x"FD", x"FC", x"00", x"04", x"02", x"FE", x"FC", x"FD", x"00", x"02", x"01",
	x"FF", x"FE", x"FB", x"F9", x"FA", x"FC", x"FC", x"FC", x"FB", x"F8", x"F5", x"F8",
	x"FE", x"02", x"00", x"FC", x"FA", x"F9", x"F9", x"FA", x"FA", x"FB", x"FE", x"01",
	x"02", x"03", x"01", x"FF", x"FD", x"FF", x"00", x"FF", x"FE", x"00", x"02", x"04",
	x"05", x"05", x"08", x"0B", x"07", x"04", x"03", x"04", x"06", x"08", x"0A", x"0C",
	x"0E", x"0E", x"0D", x"0A", x"07", x"08", x"0B", x"0C", x"0B", x"0A", x"0A", x"08",
	x"05", x"03", x"06", x"0B", x"0D", x"0A", x"08", x"08", x"08", x"04", x"00", x"01",
	x"05", x"07", x"05", x"02", x"01", x"03", x"04", x"01", x"FC", x"FA", x"F9", x"F6",
	x"F5", x"F7", x"F8", x"F8", x"F9", x"F7", x"F4", x"F8", x"FD", x"FC", x"FB", x"FB",
	x"FB", x"F9", x"F8", x"F9", x"FB", x"FD", x"FE", x"FD", x"FE", x"00", x"FF", x"00",
	x"03", x"06", x"05", x"01", x"FE", x"FB", x"F9", x"F8", x"F9", x"FD", x"FF", x"FF",
	x"01", x"02", x"FF", x"FD", x"FD", x"FE", x"FE", x"FD", x"FE", x"01", x"04", x"05",
	x"03", x"01", x"FE", x"FC", x"FB", x"FB", x"FA", x"F7", x"F5", x"F3", x"F3", x"F5",
	x"F7", x"F6", x"F7", x"F9", x"F8", x"F7", x"F7", x"F8", x"FB", x"FB", x"F9", x"FA",
	x"FB", x"FD", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"FB", x"FA", x"FE", x"02",
	x"02", x"01", x"00", x"01", x"03", x"04", x"05", x"04", x"02", x"01", x"01", x"02",
	x"04", x"07", x"0B", x"0B", x"06", x"00", x"FE", x"FF", x"01", x"00", x"FE", x"FC",
	x"F9", x"F9", x"FB", x"FE", x"00", x"01", x"00", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"02", x"05", x"05", x"02", x"00", x"01", x"03", x"04", x"04", x"04", x"03",
	x"04", x"05", x"04", x"01", x"00", x"00", x"03", x"05", x"06", x"05", x"05", x"07",
	x"06", x"03", x"01", x"FF", x"FF", x"00", x"01", x"02", x"02", x"02", x"01", x"00",
	x"00", x"FE", x"FD", x"FF", x"01", x"01", x"02", x"03", x"01", x"FD", x"FA", x"FA",
	x"FD", x"01", x"02", x"FE", x"FA", x"F8", x"FA", x"FC", x"F9", x"F8", x"FB", x"FE",
	x"FC", x"FB", x"FB", x"FC", x"FC", x"FC", x"FA", x"F8", x"F9", x"FD", x"02", x"03",
	x"00", x"FC", x"FB", x"FE", x"00", x"00", x"00", x"01", x"FE", x"FB", x"FC", x"01",
	x"01", x"FD", x"FD", x"01", x"06", x"06", x"04", x"03", x"02", x"01", x"01", x"03",
	x"03", x"00", x"FD", x"FE", x"FF", x"FE", x"FE", x"00", x"FF", x"FA", x"F9", x"FC",
	x"FC", x"F9", x"F9", x"FB", x"FA", x"FA", x"FD", x"FE", x"FD", x"FD", x"FF", x"FF",
	x"FE", x"FD", x"00", x"05", x"05", x"03", x"03", x"04", x"05", x"06", x"05", x"02",
	x"FE", x"FD", x"00", x"02", x"00", x"01", x"04", x"05", x"02", x"FD", x"FA", x"FC",
	x"00", x"04", x"06", x"06", x"05", x"04", x"04", x"04", x"03", x"00", x"FF", x"01",
	x"02", x"00", x"FD", x"FD", x"01", x"02", x"01", x"03", x"06", x"08", x"07", x"05",
	x"04", x"05", x"03", x"03", x"04", x"03", x"01", x"FF", x"FE", x"FE", x"02", x"04",
	x"FF", x"F8", x"F6", x"FA", x"FC", x"F9", x"F6", x"F6", x"F9", x"FB", x"FC", x"FB",
	x"FA", x"FB", x"FB", x"FD", x"FE", x"FF", x"FF", x"FE", x"FD", x"FC", x"FB", x"FA",
	x"F9", x"F8", x"FA", x"FC", x"FD", x"FB", x"FB", x"FE", x"FF", x"FD", x"FC", x"FC",
	x"FC", x"FD", x"FE", x"FF", x"00", x"01", x"00", x"FF", x"FF", x"00", x"02", x"04",
	x"02", x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"FF", x"FB", x"F8", x"F8", x"FA",
	x"FD", x"FD", x"FB", x"F9", x"F6", x"F5", x"F6", x"FB", x"FF", x"00", x"00", x"00",
	x"FD", x"FD", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FD", x"FF", x"01",
	x"02", x"02", x"02", x"04", x"07", x"04", x"FF", x"FF", x"03", x"04", x"00", x"FF",
	x"03", x"05", x"04", x"02", x"02", x"05", x"06", x"04", x"01", x"FE", x"00", x"02",
	x"04", x"05", x"04", x"03", x"02", x"01", x"01", x"01", x"03", x"03", x"01", x"02",
	x"04", x"04", x"04", x"06", x"0A", x"0C", x"0B", x"09", x"07", x"07", x"08", x"07",
	x"06", x"09", x"0C", x"0A", x"08", x"06", x"04", x"01", x"FE", x"FC", x"FD", x"FE",
	x"00", x"00", x"FF", x"FC", x"FA", x"FA", x"FB", x"F8", x"F6", x"FA", x"FE", x"FC",
	x"F9", x"FC", x"FF", x"FD", x"FB", x"FC", x"FD", x"FB", x"FA", x"FB", x"FB", x"FA",
	x"F9", x"FB", x"FE", x"FF", x"00", x"FF", x"FE", x"FE", x"FF", x"02", x"05", x"06",
	x"05", x"02", x"FD", x"FA", x"FB", x"FC", x"FC", x"FC", x"FE", x"FF", x"00", x"01",
	x"FF", x"FF", x"FD", x"FA", x"F8", x"F9", x"F9", x"F9", x"FB", x"FD", x"FD", x"FB",
	x"FB", x"FC", x"FB", x"FB", x"FC", x"FB", x"FB", x"FB", x"FB", x"FC", x"FE", x"FE",
	x"FB", x"F9", x"FB", x"FF", x"00", x"FD", x"FA", x"F9", x"FA", x"FA", x"FB", x"00",
	x"04", x"05", x"02", x"02", x"05", x"07", x"04", x"02", x"04", x"08", x"08", x"04",
	x"FF", x"FF", x"02", x"01", x"FD", x"FD", x"00", x"04", x"03", x"01", x"01", x"04",
	x"08", x"07", x"03", x"02", x"02", x"00", x"00", x"02", x"05", x"03", x"FE", x"FB",
	x"FB", x"FB", x"FB", x"FB", x"FB", x"F7", x"F3", x"F1", x"F2", x"F6", x"F8", x"F8",
	x"F9", x"F9", x"FB", x"FE", x"01", x"05", x"07", x"04", x"02", x"02", x"04", x"07",
	x"06", x"02", x"02", x"04", x"04", x"03", x"03", x"04", x"03", x"01", x"FF", x"00",
	x"03", x"02", x"FD", x"FC", x"FF", x"02", x"04", x"05", x"05", x"04", x"02", x"01",
	x"00", x"00", x"01", x"02", x"02", x"02", x"01", x"00", x"FF", x"FE", x"FE", x"FD",
	x"FB", x"FB", x"FC", x"FB", x"FB", x"FD", x"FD", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FC", x"FF", x"01", x"FF", x"FE", x"FE", x"FC", x"FB", x"FD", x"00", x"FE", x"FB",
	x"FC", x"01", x"04", x"00", x"FD", x"FE", x"00", x"00", x"FE", x"FE", x"FE", x"00",
	x"01", x"00", x"FE", x"FC", x"FF", x"03", x"04", x"03", x"01", x"02", x"02", x"02",
	x"03", x"04", x"02", x"01", x"02", x"04", x"04", x"04", x"01", x"FD", x"FA", x"FB",
	x"FD", x"FE", x"FC", x"FB", x"FB", x"FC", x"FD", x"FE", x"00", x"00", x"FE", x"FE",
	x"01", x"02", x"FF", x"FC", x"FB", x"FB", x"FB", x"F9", x"F8", x"F9", x"FE", x"02",
	x"03", x"00", x"FD", x"FD", x"FE", x"00", x"01", x"02", x"03", x"04", x"08", x"0D",
	x"0E", x"0E", x"0E", x"0F", x"0E", x"0A", x"07", x"07", x"06", x"06", x"05", x"04",
	x"04", x"06", x"07", x"05", x"04", x"06", x"06", x"05", x"02", x"FF", x"FE", x"FD",
	x"FC", x"FC", x"FD", x"FD", x"FB", x"F9", x"F8", x"F9", x"F9", x"F9", x"F9", x"F8",
	x"F7", x"F7", x"F8", x"FB", x"FA", x"F5", x"F2", x"F3", x"F7", x"FC", x"FE", x"FE",
	x"00", x"02", x"00", x"FB", x"FA", x"FF", x"03", x"02", x"FF", x"FE", x"FE", x"FF",
	x"02", x"03", x"00", x"FF", x"00", x"00", x"FE", x"FC", x"FC", x"FC", x"FC", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"00", x"FE", x"FC", x"FC", x"FE", x"FD", x"FB", x"FC",
	x"00", x"04", x"04", x"00", x"FC", x"FC", x"FC", x"FA", x"FA", x"FB", x"FE", x"00",
	x"FD", x"F7", x"F4", x"F6", x"F9", x"FC", x"FE", x"FE", x"FF", x"FF", x"FE", x"FB",
	x"F9", x"FB", x"FF", x"01", x"FF", x"FD", x"FE", x"02", x"06", x"04", x"00", x"FF",
	x"02", x"05", x"06", x"06", x"06", x"06", x"06", x"07", x"08", x"08", x"07", x"07",
	x"06", x"04", x"02", x"02", x"06", x"08", x"07", x"05", x"05", x"04", x"02", x"01",
	x"02", x"02", x"00", x"FE", x"FC", x"F9", x"F6", x"F8", x"FB", x"FB", x"FB", x"FA",
	x"FC", x"FF", x"FE", x"FC", x"FE", x"01", x"00", x"FE", x"FB", x"FA", x"FD", x"00",
	x"02", x"04", x"05", x"06", x"06", x"04", x"01", x"01", x"02", x"01", x"01", x"02",
	x"04", x"05", x"04", x"03", x"04", x"05", x"04", x"03", x"01", x"FF", x"FE", x"FE",
	x"00", x"03", x"03", x"02", x"02", x"01", x"FF", x"00", x"05", x"07", x"04", x"00",
	x"FF", x"00", x"FE", x"FB", x"FC", x"FF", x"02", x"01", x"FF", x"FE", x"FD", x"FA",
	x"F7", x"F6", x"F6", x"F5", x"F4", x"F7", x"FA", x"FB", x"FB", x"FB", x"FA", x"F8",
	x"F8", x"F7", x"F6", x"F8", x"FB", x"FF", x"00", x"FE", x"FC", x"FC", x"FD", x"FD",
	x"FC", x"FD", x"FF", x"FF", x"00", x"03", x"05", x"04", x"00", x"FF", x"01", x"03",
	x"03", x"04", x"04", x"06", x"07", x"05", x"04", x"05", x"08", x"0A", x"06", x"01",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FB", x"F9", x"F9", x"F9", x"FC", x"FF",
	x"FF", x"FB", x"F8", x"F9", x"FB", x"FD", x"01", x"02", x"00", x"FE", x"FF", x"FF",
	x"FF", x"01", x"01", x"FF", x"FB", x"F9", x"FB", x"FF", x"02", x"03", x"03", x"04",
	x"05", x"05", x"02", x"02", x"03", x"02", x"FF", x"FD", x"FF", x"03", x"04", x"04",
	x"04", x"04", x"03", x"02", x"02", x"03", x"03", x"03", x"01", x"FD", x"FD", x"FF",
	x"04", x"05", x"03", x"04", x"03", x"00", x"FE", x"01", x"02", x"01", x"FF", x"FE",
	x"FE", x"FC", x"F9", x"FA", x"FB", x"FA", x"F7", x"F6", x"F7", x"F6", x"F8", x"FC",
	x"00", x"03", x"01", x"FD", x"FC", x"FE", x"00", x"FD", x"F9", x"FA", x"FE", x"02",
	x"01", x"FE", x"FD", x"FD", x"FE", x"00", x"02", x"00", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"00", x"01", x"02", x"02", x"01", x"01", x"03", x"02", x"FF", x"FE", x"00",
	x"00", x"FE", x"FF", x"03", x"06", x"07", x"03", x"01", x"00", x"FF", x"FF", x"00",
	x"FF", x"01", x"02", x"01", x"FF", x"FC", x"FE", x"00", x"01", x"02", x"03", x"04",
	x"02", x"FF", x"FE", x"FF", x"00", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF",
	x"00", x"FF", x"FC", x"FC", x"FD", x"FD", x"FD", x"FE", x"00", x"01", x"02", x"02",
	x"02", x"01", x"00", x"FF", x"FF", x"01", x"03", x"04", x"04", x"04", x"05", x"02",
	x"FE", x"FF", x"02", x"01", x"FF", x"FF", x"02", x"03", x"00", x"FB", x"FB", x"FD",
	x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FF", x"02", x"02", x"01", x"00", x"00",
	x"00", x"FE", x"FC", x"FE", x"00", x"01", x"02", x"04", x"06", x"05", x"02", x"01",
	x"00", x"FF", x"FD", x"FA", x"F9", x"FA", x"FB", x"FD", x"FF", x"02", x"03", x"04",
	x"03", x"01", x"FD", x"FD", x"FE", x"FE", x"FD", x"FD", x"FC", x"FD", x"00", x"01",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FD", x"FC",
	x"FC", x"FE", x"FF", x"FE", x"FE", x"FF", x"01", x"02", x"02", x"02", x"00", x"FD",
	x"FB", x"FB", x"FA", x"F7", x"F9", x"FD", x"FE", x"FB", x"F8", x"F6", x"F6", x"F7",
	x"F7", x"F8", x"F8", x"F8", x"FA", x"FF", x"01", x"FE", x"FD", x"02", x"05", x"04",
	x"02", x"03", x"03", x"02", x"FF", x"00", x"05", x"07", x"07", x"05", x"04", x"03",
	x"02", x"02", x"03", x"03", x"01", x"FF", x"02", x"05", x"05", x"03", x"02", x"04",
	x"06", x"04", x"03", x"01", x"FF", x"FD", x"FD", x"FE", x"FF", x"FF", x"01", x"03",
	x"05", x"04", x"02", x"02", x"02", x"FF", x"FB", x"FB", x"00", x"02", x"01", x"00",
	x"FF", x"FF", x"00", x"02", x"03", x"03", x"02", x"00", x"FE", x"FD", x"FE", x"FE",
	x"FF", x"FE", x"FB", x"FB", x"FD", x"FF", x"FF", x"FF", x"FE", x"FD", x"FC", x"FD",
	x"FF", x"02", x"03", x"02", x"00", x"00", x"00", x"FE", x"FE", x"00", x"01", x"FF",
	x"FE", x"00", x"03", x"05", x"04", x"01", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"01", x"00", x"FD", x"FB", x"FD", x"FB", x"F8", x"F7", x"FB", x"FD", x"FC", x"F9",
	x"F8", x"F9", x"F8", x"F7", x"FB", x"01", x"03", x"FF", x"F9", x"F6", x"F7", x"F9",
	x"FC", x"FE", x"FF", x"FC", x"FA", x"FA", x"FE", x"03", x"02", x"FF", x"FF", x"03",
	x"02", x"FF", x"01", x"02", x"02", x"01", x"01", x"01", x"03", x"06", x"07", x"07",
	x"06", x"05", x"05", x"06", x"07", x"07", x"06", x"04", x"03", x"03", x"05", x"06",
	x"05", x"01", x"FE", x"FE", x"FF", x"FE", x"FD", x"FD", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FC", x"FB", x"FC", x"FC", x"F9", x"F8", x"FA", x"F9", x"F5", x"F4",
	x"F9", x"FF", x"02", x"01", x"FE", x"FD", x"FD", x"FB", x"FB", x"FE", x"00", x"00",
	x"00", x"FF", x"00", x"01", x"FF", x"FE", x"FF", x"01", x"01", x"01", x"00", x"01",
	x"01", x"00", x"FE", x"FE", x"00", x"05", x"08", x"06", x"03", x"03", x"03", x"04",
	x"03", x"02", x"02", x"03", x"01", x"00", x"01", x"03", x"04", x"05", x"04", x"00",
	x"FD", x"FB", x"FF", x"04", x"05", x"02", x"00", x"FF", x"FC", x"FA", x"F9", x"F8",
	x"F8", x"F8", x"F8", x"F8", x"F8", x"F9", x"F9", x"FA", x"FB", x"FC", x"FA", x"FA",
	x"FE", x"00", x"FF", x"FE", x"FE", x"00", x"02", x"02", x"03", x"04", x"03", x"02",
	x"03", x"04", x"03", x"02", x"03", x"08", x"0A", x"05", x"01", x"00", x"00", x"FD",
	x"FA", x"FB", x"FC", x"FC", x"FB", x"FA", x"FA", x"FD", x"FF", x"FD", x"FA", x"FB",
	x"FD", x"FE", x"FB", x"FB", x"FF", x"00", x"FE", x"FE", x"FF", x"FF", x"FE", x"FD",
	x"FC", x"FD", x"00", x"00", x"FF", x"FF", x"FE", x"FD", x"FE", x"FE", x"FE", x"00",
	x"01", x"00", x"FC", x"FC", x"01", x"04", x"04", x"00", x"FF", x"01", x"02", x"03",
	x"03", x"03", x"02", x"01", x"03", x"05", x"06", x"06", x"08", x"0A", x"08", x"05",
	x"05", x"07", x"09", x"08", x"06", x"04", x"04", x"04", x"04", x"02", x"04", x"04",
	x"05", x"05", x"01", x"FA", x"F8", x"FC", x"01", x"03", x"00", x"FE", x"00", x"01",
	x"FD", x"F6", x"F4", x"F6", x"F9", x"F8", x"F4", x"F3", x"F9", x"FE", x"FF", x"FD",
	x"FD", x"FD", x"FC", x"FC", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"02", x"03", x"02", x"01", x"01", x"02", x"05", x"05",
	x"03", x"01", x"FF", x"FE", x"FE", x"FE", x"FF", x"02", x"02", x"FF", x"FE", x"FE",
	x"FC", x"FC", x"FE", x"FF", x"FE", x"FC", x"FE", x"02", x"03", x"00", x"FE", x"FE",
	x"FC", x"F9", x"F6", x"F4", x"F3", x"F6", x"FA", x"FD", x"FD", x"FD", x"FC", x"FB",
	x"FC", x"01", x"04", x"02", x"FE", x"FC", x"FC", x"FD", x"FE", x"00", x"03", x"05",
	x"04", x"03", x"03", x"02", x"01", x"01", x"03", x"05", x"07", x"07", x"07", x"09",
	x"0A", x"09", x"05", x"03", x"04", x"02", x"FE", x"FF", x"01", x"00", x"FE", x"FF",
	x"01", x"00", x"FC", x"F7", x"F8", x"FB", x"FE", x"FF", x"FD", x"FB", x"FB", x"FA",
	x"FA", x"FA", x"FA", x"FA", x"FB", x"FA", x"FB", x"FB", x"FC", x"FE", x"FE", x"FC",
	x"FB", x"FD", x"FE", x"FE", x"FE", x"00", x"03", x"01", x"FC", x"FB", x"FE", x"FF",
	x"FD", x"FD", x"00", x"04", x"04", x"03", x"04", x"06", x"06", x"04", x"03", x"04",
	x"04", x"03", x"03", x"03", x"02", x"01", x"04", x"06", x"03", x"00", x"FF", x"FF",
	x"FE", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"FC", x"F9", x"FB", x"FE", x"FE",
	x"FB", x"FB", x"FD", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"01",
	x"02", x"00", x"FE", x"FF", x"04", x"05", x"04", x"02", x"02", x"01", x"FF", x"FE",
	x"FF", x"FF", x"00", x"FF", x"FC", x"FB", x"FB", x"FC", x"FD", x"FF", x"FE", x"FC",
	x"FC", x"00", x"03", x"03", x"02", x"03", x"03", x"01", x"00", x"01", x"02", x"01",
	x"FF", x"FC", x"F9", x"F9", x"FB", x"FC", x"FC", x"F9", x"F9", x"FC", x"FB", x"F7",
	x"F7", x"FA", x"FD", x"FC", x"FB", x"FC", x"00", x"02", x"01", x"FF", x"FD", x"FE",
	x"00", x"02", x"03", x"04", x"04", x"05", x"05", x"05", x"05", x"05", x"04", x"05",
	x"05", x"03", x"01", x"01", x"03", x"05", x"04", x"03", x"01", x"00", x"01", x"03",
	x"04", x"04", x"01", x"00", x"00", x"02", x"04", x"04", x"05", x"05", x"02", x"FE",
	x"FC", x"FD", x"FF", x"00", x"FF", x"FD", x"FB", x"FA", x"F9", x"F8", x"F9", x"FD",
	x"FF", x"FE", x"FC", x"FA", x"F7", x"F7", x"FB", x"FE", x"FE", x"FC", x"FA", x"FB",
	x"FE", x"FF", x"00", x"02", x"05", x"06", x"05", x"03", x"03", x"04", x"03", x"02",
	x"02", x"02", x"01", x"01", x"01", x"02", x"00", x"FF", x"FD", x"FA", x"FB", x"FC",
	x"FD", x"FC", x"FC", x"FD", x"00", x"03", x"02", x"FC", x"F7", x"F9", x"FC", x"FD",
	x"FC", x"FB", x"FC", x"FB", x"FA", x"F9", x"FA", x"FE", x"FF", x"FD", x"FC", x"FE",
	x"01", x"02", x"01", x"FF", x"FF", x"FF", x"FE", x"FD", x"FF", x"02", x"04", x"03",
	x"01", x"02", x"03", x"03", x"00", x"FD", x"FE", x"01", x"02", x"00", x"FE", x"00",
	x"02", x"01", x"02", x"03", x"05", x"05", x"05", x"02", x"FF", x"FD", x"FC", x"FE",
	x"00", x"01", x"00", x"00", x"01", x"01", x"01", x"00", x"01", x"03", x"02", x"01",
	x"FF", x"FE", x"FC", x"FC", x"FC", x"FB", x"FB", x"FD", x"FC", x"FB", x"FE", x"00",
	x"FE", x"FC", x"F9", x"F9", x"FA", x"FA", x"FB", x"FD", x"FE", x"FE", x"FE", x"FE",
	x"00", x"01", x"01", x"01", x"01", x"01", x"FF", x"00", x"02", x"03", x"01", x"00",
	x"00", x"01", x"01", x"02", x"01", x"02", x"04", x"05", x"04", x"05", x"04", x"01",
	x"FF", x"01", x"04", x"03", x"01", x"04", x"05", x"03", x"01", x"01", x"03", x"04",
	x"04", x"04", x"06", x"07", x"06", x"04", x"06", x"07", x"05", x"01", x"00", x"01",
	x"FF", x"FD", x"FC", x"FB", x"FA", x"F9", x"FB", x"FE", x"00", x"FD", x"FB", x"FB",
	x"FB", x"FB", x"FB", x"FA", x"F8", x"F9", x"FC", x"FB", x"FA", x"F9", x"FB", x"FB",
	x"F9", x"F8", x"FA", x"FB", x"F9", x"F9", x"FD", x"00", x"00", x"02", x"05", x"04",
	x"FD", x"F7", x"F9", x"FF", x"02", x"02", x"01", x"FF", x"FE", x"FF", x"01", x"01",
	x"FF", x"FE", x"FD", x"FB", x"FB", x"FC", x"FF", x"00", x"FF", x"00", x"00", x"FC",
	x"FC", x"01", x"02", x"FE", x"F9", x"F8", x"FB", x"FE", x"FF", x"00", x"02", x"03",
	x"01", x"00", x"03", x"06", x"04", x"FF", x"FD", x"FD", x"FD", x"FD", x"FC", x"FD",
	x"FE", x"FE", x"FD", x"FF", x"04", x"06", x"04", x"00", x"FF", x"FF", x"01", x"02",
	x"03", x"02", x"01", x"01", x"02", x"04", x"04", x"04", x"03", x"01", x"01", x"03",
	x"05", x"04", x"03", x"03", x"00", x"FB", x"F8", x"FA", x"FD", x"FF", x"01", x"03",
	x"03", x"02", x"00", x"FF", x"FF", x"FD", x"FB", x"FE", x"FF", x"FE", x"FF", x"00",
	x"00", x"FF", x"03", x"06", x"04", x"01", x"01", x"02", x"01", x"00", x"FF", x"FF",
	x"FD", x"FB", x"FB", x"FF", x"01", x"00", x"FF", x"FF", x"FD", x"F8", x"F7", x"F8",
	x"F9", x"F9", x"FB", x"FD", x"FD", x"FF", x"01", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"00", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"04", x"06",
	x"06", x"08", x"0A", x"07", x"01", x"00", x"01", x"01", x"02", x"01", x"01", x"01",
	x"02", x"00", x"FF", x"FD", x"FC", x"FC", x"FC", x"FB", x"FB", x"FC", x"FD", x"FB",
	x"FB", x"FC", x"FD", x"FD", x"FC", x"FF", x"01", x"00", x"FF", x"FF", x"00", x"00",
	x"FE", x"FD", x"FC", x"FC", x"FC", x"FC", x"FC", x"FD", x"FE", x"FF", x"FD", x"FB",
	x"FD", x"00", x"03", x"04", x"03", x"01", x"FF", x"00", x"05", x"06", x"01", x"FC",
	x"FC", x"FE", x"FF", x"00", x"01", x"01", x"01", x"00", x"FE", x"FC", x"FC", x"FE",
	x"00", x"02", x"03", x"01", x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"FF", x"FD",
	x"FD", x"FE", x"00", x"FF", x"FC", x"FC", x"FC", x"FB", x"FA", x"FB", x"FE", x"01",
	x"01", x"03", x"03", x"02", x"01", x"02", x"02", x"03", x"03", x"03", x"04", x"02",
	x"01", x"02", x"07", x"0B", x"0C", x"0B", x"0A", x"08", x"05", x"02", x"01", x"FF",
	x"FD", x"FC", x"FC", x"FD", x"FD", x"FC", x"FE", x"00", x"00", x"FD", x"FA", x"F8",
	x"F8", x"F9", x"FA", x"FD", x"01", x"00", x"FC", x"FD", x"FF", x"FD", x"F9", x"F8",
	x"FA", x"FB", x"FB", x"FA", x"F8", x"F5", x"F5", x"F7", x"FA", x"FB", x"FB", x"FD",
	x"FF", x"FE", x"FB", x"FA", x"FB", x"FD", x"FB", x"FB", x"FD", x"00", x"00", x"00",
	x"02", x"03", x"02", x"02", x"03", x"03", x"04", x"05", x"03", x"01", x"01", x"03",
	x"04", x"04", x"03", x"02", x"03", x"05", x"07", x"07", x"06", x"05", x"04", x"02",
	x"02", x"02", x"04", x"03", x"02", x"01", x"01", x"01", x"01", x"01", x"00", x"FC",
	x"FA", x"FC", x"FF", x"01", x"00", x"FE", x"FB", x"FA", x"FB", x"FF", x"02", x"01",
	x"FF", x"00", x"03", x"02", x"FF", x"FD", x"00", x"FF", x"FA", x"F7", x"F8", x"FA",
	x"FE", x"01", x"FE", x"FC", x"FD", x"FE", x"00", x"03", x"04", x"04", x"01", x"00",
	x"03", x"05", x"05", x"04", x"06", x"08", x"04", x"00", x"00", x"03", x"05", x"04",
	x"00", x"FD", x"FD", x"FD", x"FC", x"FD", x"FE", x"FC", x"FC", x"FD", x"FE", x"FE",
	x"FD", x"F9", x"F8", x"FB", x"FE", x"FD", x"FC", x"FB", x"FC", x"FC", x"FA", x"F8",
	x"F8", x"FB", x"FB", x"F7", x"F5", x"F5", x"F6", x"F7", x"F9", x"FB", x"FD", x"FE",
	x"01", x"03", x"04", x"05", x"05", x"05", x"08", x"0A", x"0A", x"09", x"08", x"06",
	x"04", x"01", x"03", x"06", x"06", x"03", x"00", x"FF", x"FE", x"FD", x"FD", x"FE",
	x"FE", x"FD", x"00", x"03", x"01", x"FE", x"FE", x"FD", x"FB", x"FB", x"FD", x"FF",
	x"00", x"01", x"01", x"00", x"FE", x"FD", x"FC", x"FC", x"FC", x"FB", x"FA", x"FB",
	x"FD", x"FE", x"FE", x"FF", x"00", x"FE", x"FD", x"FE", x"00", x"00", x"FE", x"FD",
	x"FE", x"01", x"FF", x"FC", x"FD", x"00", x"03", x"01", x"FE", x"FD", x"00", x"04",
	x"04", x"02", x"00", x"FF", x"FF", x"00", x"01", x"01", x"01", x"03", x"05", x"05",
	x"05", x"08", x"0A", x"06", x"03", x"01", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FC", x"FB", x"FC", x"FE", x"FE",
	x"FE", x"00", x"03", x"05", x"06", x"06", x"09", x"09", x"07", x"05", x"04", x"03",
	x"01", x"00", x"01", x"05", x"06", x"04", x"02", x"01", x"01", x"01", x"00", x"FF",
	x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FD", x"FE", x"01", x"03", x"00", x"FE",
	x"FF", x"01", x"FF", x"FC", x"FB", x"FC", x"FD", x"FE", x"FB", x"FA", x"FA", x"F9",
	x"F7", x"F7", x"FA", x"FD", x"FD", x"FB", x"F9", x"F7", x"F6", x"F8", x"F8", x"F7",
	x"F7", x"F7", x"F5", x"F3", x"F5", x"F9", x"FB", x"F9", x"FA", x"FC", x"FC", x"FA",
	x"FA", x"FD", x"FF", x"FE", x"FB", x"FB", x"FC", x"FD", x"FF", x"02", x"04", x"05",
	x"06", x"08", x"09", x"08", x"07", x"07", x"06", x"05", x"04", x"04", x"04", x"07",
	x"09", x"08", x"05", x"05", x"05", x"05", x"04", x"03", x"02", x"02", x"00", x"FF",
	x"FF", x"00", x"FF", x"FE", x"FE", x"00", x"02", x"01", x"FD", x"FB", x"FA", x"FA",
	x"FB", x"FB", x"FB", x"FB", x"FC", x"FD", x"FC", x"FD", x"00", x"01", x"FE", x"FB",
	x"FC", x"FD", x"FD", x"FD", x"00", x"03", x"02", x"FF", x"FD", x"FD", x"FD", x"FC",
	x"FD", x"00", x"01", x"02", x"02", x"04", x"05", x"04", x"02", x"03", x"05", x"04",
	x"03", x"04", x"05", x"04", x"03", x"00", x"FC", x"FA", x"FD", x"FF", x"FE", x"FC",
	x"FD", x"FE", x"FC", x"FA", x"FA", x"FC", x"FD", x"FB", x"FA", x"FA", x"FD", x"FF",
	x"FC", x"FC", x"FE", x"FF", x"FE", x"FC", x"FC", x"FE", x"00", x"02", x"03", x"02",
	x"FE", x"FA", x"FB", x"00", x"03", x"03", x"03", x"03", x"04", x"04", x"04", x"04",
	x"07", x"09", x"09", x"07", x"05", x"04", x"03", x"04", x"05", x"05", x"04", x"03",
	x"01", x"FD", x"FC", x"FE", x"FE", x"FC", x"F9", x"F9", x"F9", x"F8", x"F6", x"F7",
	x"F9", x"FB", x"FD", x"FF", x"01", x"03", x"04", x"02", x"FF", x"FD", x"FD", x"FE",
	x"FE", x"FD", x"FD", x"FF", x"00", x"01", x"FF", x"FE", x"FE", x"FC", x"FB", x"FC",
	x"FC", x"FC", x"FA", x"FA", x"FB", x"FE", x"FE", x"FB", x"F9", x"F9", x"FA", x"FB",
	x"FD", x"FE", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"00", x"FF", x"00", x"02", x"03", x"02", x"01", x"02", x"03", x"03", x"00",
	x"FE", x"FE", x"00", x"03", x"04", x"05", x"05", x"05", x"03", x"03", x"04", x"05",
	x"03", x"02", x"03", x"05", x"03", x"02", x"05", x"08", x"0A", x"0A", x"08", x"05",
	x"02", x"FF", x"FD", x"FD", x"FE", x"FE", x"FF", x"FE", x"FE", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FF", x"FF", x"FD", x"FC", x"FC", x"FD",
	x"FD", x"FE", x"FD", x"FC", x"FC", x"FB", x"F8", x"F8", x"FB", x"FE", x"FF", x"FD",
	x"FB", x"FA", x"FA", x"FB", x"FD", x"FF", x"FE", x"FC", x"FC", x"FD", x"FE", x"FE",
	x"FC", x"FA", x"FA", x"FB", x"FD", x"FE", x"FE", x"00", x"00", x"00", x"FE", x"FE",
	x"FF", x"02", x"02", x"02", x"03", x"02", x"FF", x"FC", x"FD", x"FF", x"00", x"FF",
	x"00", x"02", x"04", x"06", x"07", x"06", x"04", x"01", x"02", x"05", x"06", x"05",
	x"03", x"03", x"04", x"04", x"03", x"02", x"02", x"02", x"00", x"00", x"00", x"01",
	x"01", x"02", x"02", x"FF", x"FD", x"FD", x"FF", x"01", x"01", x"00", x"01", x"02",
	x"01", x"FD", x"FB", x"FC", x"FD", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF",
	x"FD", x"FC", x"FD", x"FD", x"FD", x"FE", x"FF", x"FE", x"FE", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"01", x"01", x"FE", x"FC", x"FF", x"00", x"00",
	x"00", x"02", x"03", x"02", x"FE", x"FD", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD",
	x"FE", x"FD", x"FA", x"FA", x"FB", x"FC", x"FD", x"FD", x"FC", x"FC", x"FD", x"FF",
	x"01", x"02", x"03", x"03", x"02", x"FF", x"FE", x"00", x"03", x"04", x"01", x"FF",
	x"FE", x"FE", x"FD", x"FD", x"FD", x"FF", x"01", x"02", x"00", x"FD", x"FB", x"FB",
	x"FC", x"FE", x"01", x"03", x"04", x"02", x"01", x"00", x"FC", x"FA", x"FC", x"01",
	x"02", x"00", x"FD", x"FA", x"FA", x"FC", x"FD", x"FC", x"FC", x"FC", x"FC", x"FE",
	x"01", x"02", x"01", x"01", x"01", x"00", x"FE", x"FE", x"01", x"05", x"06", x"04",
	x"04", x"05", x"05", x"02", x"00", x"02", x"02", x"FE", x"FA", x"FA", x"FF", x"03",
	x"02", x"FD", x"FB", x"FA", x"F9", x"F8", x"FA", x"FD", x"FE", x"FE", x"FD", x"FD",
	x"FE", x"FF", x"FE", x"FD", x"FD", x"FE", x"FD", x"FA", x"FA", x"FE", x"03", x"01",
	x"FE", x"00", x"02", x"01", x"00", x"02", x"02", x"01", x"01", x"03", x"05", x"06",
	x"06", x"05", x"05", x"05", x"07", x"09", x"08", x"05", x"03", x"03", x"04", x"05",
	x"06", x"06", x"06", x"05", x"04", x"03", x"02", x"02", x"04", x"05", x"06", x"04",
	x"03", x"04", x"05", x"04", x"02", x"01", x"FE", x"FC", x"FC", x"FD", x"FE", x"00",
	x"00", x"FD", x"FA", x"FA", x"FA", x"FA", x"FB", x"FD", x"FE", x"FB", x"F9", x"FA",
	x"FD", x"FC", x"FB", x"FB", x"F9", x"F8", x"F8", x"F7", x"F8", x"FB", x"FC", x"F9",
	x"F6", x"F5", x"F8", x"FB", x"FC", x"FD", x"FD", x"FE", x"FF", x"00", x"01", x"03",
	x"02", x"01", x"01", x"01", x"01", x"03", x"03", x"01", x"00", x"02", x"02", x"00",
	x"00", x"02", x"03", x"FF", x"FA", x"FB", x"FF", x"02", x"01", x"FF", x"FF", x"01",
	x"01", x"FE", x"FD", x"FE", x"00", x"01", x"01", x"02", x"03", x"03", x"02", x"02",
	x"01", x"00", x"FD", x"FC", x"FD", x"FE", x"FE", x"FD", x"FC", x"FD", x"FD", x"FD",
	x"FD", x"FF", x"00", x"00", x"01", x"02", x"02", x"00", x"01", x"02", x"03", x"03",
	x"02", x"01", x"00", x"FF", x"01", x"03", x"02", x"FF", x"FD", x"FC", x"FC", x"FC",
	x"FD", x"00", x"02", x"03", x"03", x"03", x"02", x"02", x"02", x"00", x"01", x"02",
	x"01", x"FF", x"FB", x"F9", x"FB", x"FE", x"FE", x"FC", x"FB", x"FD", x"FD", x"FB",
	x"F8", x"F8", x"F9", x"F9", x"F8", x"F9", x"FB", x"FD", x"FD", x"FD", x"00", x"01",
	x"01", x"00", x"FF", x"FD", x"FB", x"FE", x"01", x"00", x"FD", x"FC", x"FE", x"01",
	x"03", x"03", x"03", x"05", x"06", x"05", x"02", x"01", x"04", x"07", x"07", x"04",
	x"04", x"05", x"05", x"03", x"03", x"03", x"00", x"00", x"FF", x"FC", x"FB", x"FA",
	x"FB", x"FD", x"FD", x"FB", x"FB", x"FD", x"FE", x"FE", x"00", x"00", x"FE", x"FD",
	x"FD", x"FD", x"FD", x"FF", x"02", x"03", x"03", x"01", x"FE", x"FD", x"FD", x"FC",
	x"F9", x"FB", x"FD", x"FE", x"FF", x"02", x"03", x"02", x"02", x"01", x"FE", x"FC",
	x"FC", x"FE", x"00", x"01", x"01", x"03", x"04", x"03", x"02", x"00", x"FF", x"FD",
	x"FC", x"FD", x"FD", x"FD", x"FE", x"01", x"01", x"FD", x"FB", x"FC", x"FC", x"FC",
	x"FD", x"01", x"03", x"01", x"FC", x"FB", x"FC", x"FD", x"FD", x"FD", x"00", x"02",
	x"00", x"FD", x"FF", x"02", x"02", x"FE", x"FE", x"01", x"03", x"03", x"04", x"05",
	x"07", x"06", x"03", x"01", x"02", x"04", x"04", x"05", x"08", x"09", x"08", x"05",
	x"03", x"03", x"04", x"05", x"06", x"05", x"04", x"02", x"00", x"00", x"00", x"02",
	x"03", x"01", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"00", x"FF",
	x"FE", x"FF", x"FF", x"FE", x"FD", x"FC", x"FB", x"F9", x"F7", x"F5", x"F3", x"F4",
	x"F7", x"F9", x"F9", x"FB", x"FC", x"FB", x"F9", x"F7", x"F6", x"F5", x"F6", x"F6",
	x"F5", x"F5", x"F8", x"FA", x"FA", x"F8", x"F8", x"F9", x"FB", x"FC", x"FD", x"FD",
	x"FD", x"FD", x"FC", x"FD", x"00", x"02", x"04", x"06", x"07", x"06", x"04", x"00",
	x"FE", x"01", x"04", x"05", x"04", x"04", x"03", x"02", x"02", x"04", x"06", x"06",
	x"04", x"03", x"02", x"03", x"05", x"08", x"08", x"06", x"03", x"01", x"01", x"04",
	x"05", x"04", x"02", x"01", x"FE", x"FC", x"FC", x"FE", x"01", x"04", x"03", x"01",
	x"FF", x"FD", x"FC", x"FC", x"FC", x"FE", x"00", x"01", x"01", x"FF", x"FE", x"00",
	x"01", x"02", x"02", x"01", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"01",
	x"02", x"01", x"FF", x"FF", x"01", x"02", x"00", x"00", x"01", x"01", x"FE", x"FB",
	x"F9", x"FA", x"FA", x"FB", x"FD", x"FC", x"FB", x"FC", x"FE", x"FF", x"FE", x"FD",
	x"FB", x"FA", x"FA", x"FC", x"FE", x"FD", x"FD", x"FE", x"FE", x"FE", x"00", x"01",
	x"01", x"FF", x"FD", x"FD", x"FC", x"FA", x"F9", x"FE", x"02", x"03", x"02", x"04",
	x"04", x"03", x"02", x"03", x"03", x"01", x"FF", x"00", x"02", x"02", x"01", x"02",
	x"05", x"05", x"02", x"01", x"02", x"02", x"02", x"02", x"01", x"00", x"01", x"02",
	x"01", x"01", x"01", x"04", x"04", x"01", x"FD", x"FB", x"FB", x"FB", x"FA", x"FA",
	x"FC", x"FE", x"FF", x"00", x"FD", x"FA", x"F9", x"FA", x"FD", x"FF", x"FE", x"FD",
	x"FD", x"FD", x"FC", x"FD", x"FE", x"FE", x"FD", x"FD", x"FC", x"F9", x"F9", x"FE",
	x"01", x"01", x"00", x"FF", x"FE", x"FB", x"FB", x"FC", x"FE", x"FF", x"01", x"02",
	x"02", x"01", x"01", x"02", x"04", x"04", x"00", x"FC", x"FC", x"FD", x"FD", x"00",
	x"03", x"02", x"00", x"FE", x"FC", x"FC", x"FC", x"FD", x"FE", x"FC", x"FB", x"FB",
	x"FB", x"FB", x"FF", x"03", x"07", x"08", x"04", x"01", x"00", x"01", x"02", x"04",
	x"06", x"07", x"06", x"04", x"03", x"04", x"04", x"04", x"03", x"03", x"03", x"01",
	x"FE", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"FE", x"FD", x"FE", x"00", x"03",
	x"05", x"04", x"02", x"00", x"FE", x"FF", x"00", x"02", x"02", x"01", x"00", x"FF",
	x"01", x"02", x"01", x"00", x"01", x"02", x"01", x"FF", x"FB", x"F9", x"F9", x"FA",
	x"FA", x"FA", x"FB", x"FB", x"FA", x"FA", x"FC", x"FE", x"FC", x"F8", x"F6", x"F5",
	x"F6", x"F9", x"F9", x"F7", x"F7", x"F8", x"F8", x"F7", x"F6", x"F9", x"FC", x"FE",
	x"00", x"01", x"FF", x"FC", x"FD", x"FF", x"01", x"01", x"03", x"05", x"04", x"00",
	x"FF", x"02", x"05", x"05", x"04", x"05", x"06", x"06", x"06", x"04", x"06", x"07",
	x"05", x"02", x"00", x"00", x"02", x"04", x"04", x"04", x"04", x"04", x"03", x"03",
	x"04", x"04", x"04", x"03", x"03", x"01", x"FF", x"00", x"03", x"05", x"05", x"02",
	x"00", x"FD", x"FC", x"FE", x"01", x"03", x"02", x"01", x"FF", x"FE", x"FD", x"FF",
	x"02", x"02", x"00", x"FF", x"FD", x"FC", x"FA", x"FB", x"FE", x"00", x"01", x"03",
	x"04", x"03", x"01", x"FF", x"FF", x"FE", x"FC", x"FB", x"FC", x"FE", x"FF", x"00",
	x"00", x"FF", x"FE", x"00", x"02", x"02", x"00", x"FD", x"FB", x"FB", x"FB", x"FD",
	x"FF", x"FE", x"FC", x"FE", x"00", x"01", x"00", x"00", x"01", x"00", x"FE", x"FD",
	x"FC", x"FD", x"FE", x"FE", x"FC", x"FA", x"FB", x"FE", x"00", x"02", x"01", x"01",
	x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FF", x"FC", x"FC", x"FE", x"02", x"03",
	x"01", x"00", x"00", x"01", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"01", x"01",
	x"02", x"03", x"02", x"01", x"01", x"01", x"01", x"00", x"FF", x"FC", x"FC", x"FD",
	x"FE", x"FD", x"FF", x"01", x"01", x"FF", x"FE", x"FF", x"FF", x"FE", x"FD", x"FD",
	x"FF", x"FF", x"FE", x"FE", x"00", x"01", x"00", x"FC", x"FA", x"FA", x"FC", x"FC",
	x"FB", x"FC", x"FD", x"FC", x"FB", x"FC", x"FD", x"FE", x"FD", x"FC", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FC", x"FD", x"FD", x"FC", x"FB", x"FA", x"FD", x"00", x"02",
	x"02", x"00", x"01", x"01", x"01", x"02", x"03", x"05", x"05", x"02", x"FE", x"FE",
	x"01", x"05", x"08", x"09", x"08", x"05", x"03", x"03", x"05", x"06", x"05", x"02",
	x"01", x"01", x"00", x"01", x"01", x"02", x"03", x"04", x"03", x"01", x"03", x"05",
	x"02", x"FE", x"FE", x"FE", x"FC", x"FA", x"F9", x"FB", x"FD", x"FF", x"FE", x"FD",
	x"FC", x"FD", x"FD", x"FE", x"00", x"02", x"03", x"03", x"03", x"03", x"03", x"04",
	x"04", x"03", x"01", x"00", x"FE", x"FE", x"FE", x"FE", x"FD", x"FC", x"FD", x"FB",
	x"F7", x"F6", x"F8", x"FA", x"F8", x"F9", x"FC", x"FE", x"FB", x"F9", x"F9", x"FA",
	x"FA", x"FA", x"FB", x"FC", x"FB", x"FC", x"00", x"02", x"01", x"01", x"01", x"FF",
	x"FC", x"FB", x"FC", x"FD", x"FE", x"FF", x"02", x"05", x"02", x"FC", x"FC", x"01",
	x"04", x"03", x"02", x"01", x"00", x"00", x"03", x"06", x"06", x"05", x"04", x"02",
	x"01", x"02", x"01", x"01", x"02", x"04", x"04", x"02", x"00", x"01", x"03", x"04",
	x"05", x"04", x"02", x"FF", x"FF", x"01", x"03", x"03", x"04", x"04", x"04", x"03",
	x"03", x"03", x"02", x"02", x"02", x"01", x"FF", x"FE", x"00", x"00", x"FF", x"FF",
	x"00", x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"02", x"01", x"FF", x"FC", x"FA",
	x"F9", x"F9", x"FB", x"FC", x"FC", x"FB", x"FC", x"FD", x"FD", x"FE", x"FD", x"FC",
	x"FA", x"FA", x"FA", x"FB", x"FD", x"FE", x"FD", x"FD", x"FE", x"FD", x"FC", x"FC",
	x"FD", x"FD", x"FC", x"FD", x"FF", x"01", x"00", x"FF", x"00", x"02", x"03", x"02",
	x"02", x"03", x"03", x"04", x"04", x"04", x"03", x"02", x"02", x"02", x"01", x"01",
	x"01", x"02", x"01", x"00", x"00", x"01", x"02", x"01", x"FE", x"FD", x"FF", x"00",
	x"FF", x"FC", x"FA", x"FA", x"FA", x"FB", x"FC", x"FE", x"01", x"01", x"FE", x"FD",
	x"FF", x"01", x"02", x"01", x"01", x"01", x"00", x"FF", x"FD", x"FD", x"00", x"02",
	x"03", x"03", x"01", x"FF", x"FE", x"FE", x"FF", x"FD", x"FB", x"FB", x"FD", x"FD",
	x"FC", x"FC", x"FD", x"00", x"00", x"FE", x"FE", x"FF", x"00", x"FF", x"FD", x"FC",
	x"FE", x"00", x"00", x"FF", x"FD", x"FB", x"F9", x"F9", x"FA", x"FB", x"FA", x"FA",
	x"FB", x"FD", x"FC", x"FB", x"FB", x"FE", x"00", x"FF", x"FE", x"00", x"01", x"00",
	x"01", x"01", x"01", x"01", x"02", x"02", x"04", x"07", x"07", x"06", x"05", x"04",
	x"04", x"04", x"05", x"04", x"04", x"06", x"07", x"06", x"07", x"07", x"07", x"06",
	x"06", x"04", x"02", x"02", x"04", x"03", x"01", x"FF", x"FF", x"FE", x"FF", x"00",
	x"01", x"00", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"01", x"02",
	x"01", x"FF", x"FF", x"00", x"FF", x"FB", x"F8", x"F9", x"FC", x"FE", x"FE", x"FD",
	x"FD", x"FC", x"FC", x"FC", x"FB", x"F9", x"F9", x"FA", x"FA", x"F9", x"FA", x"FA",
	x"FB", x"FD", x"FF", x"FF", x"FF", x"00", x"00", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FD", x"FC", x"FC", x"FC", x"FD", x"FC", x"FC", x"FE", x"FF", x"00", x"FF",
	x"FE", x"FD", x"FB", x"FA", x"FC", x"00", x"01", x"00", x"00", x"01", x"02", x"02",
	x"01", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FE", x"01", x"03",
	x"03", x"02", x"03", x"03", x"01", x"FF", x"00", x"01", x"01", x"01", x"03", x"05",
	x"04", x"02", x"03", x"05", x"04", x"02", x"01", x"02", x"02", x"01", x"01", x"02",
	x"03", x"04", x"03", x"03", x"03", x"03", x"03", x"03", x"04", x"02", x"01", x"00",
	x"01", x"FF", x"FD", x"FC", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"00", x"FF",
	x"FB", x"F7", x"F4", x"F4", x"F6", x"F8", x"F9", x"FB", x"FC", x"FC", x"FC", x"FC",
	x"FC", x"FB", x"FB", x"FD", x"FC", x"FB", x"FC", x"FD", x"FD", x"FC", x"FD", x"FD",
	x"FD", x"FD", x"FC", x"FA", x"FA", x"FD", x"FF", x"FF", x"FE", x"FE", x"FF", x"00",
	x"00", x"00", x"01", x"04", x"05", x"05", x"05", x"05", x"03", x"03", x"03", x"02",
	x"03", x"05", x"06", x"04", x"02", x"02", x"02", x"02", x"02", x"04", x"05", x"04",
	x"02", x"01", x"01", x"01", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"01", x"03", x"02", x"00", x"FE", x"FC", x"FA", x"F7",
	x"F8", x"FA", x"FB", x"F9", x"F9", x"FB", x"FB", x"FB", x"FB", x"FD", x"FD", x"FC",
	x"FB", x"FC", x"FE", x"00", x"02", x"03", x"02", x"00", x"FF", x"00", x"02", x"04",
	x"04", x"04", x"02", x"02", x"03", x"02", x"00", x"FF", x"FF", x"00", x"FF", x"FE",
	x"FD", x"FC", x"FC", x"FD", x"FD", x"FE", x"FE", x"00", x"00", x"FD", x"FE", x"01",
	x"03", x"02", x"02", x"03", x"04", x"03", x"04", x"04", x"01", x"00", x"01", x"04",
	x"06", x"05", x"05", x"05", x"05", x"05", x"04", x"03", x"01", x"02", x"03", x"01",
	x"00", x"00", x"02", x"04", x"04", x"02", x"00", x"FF", x"FF", x"00", x"00", x"FF",
	x"FE", x"FE", x"FE", x"FD", x"FB", x"FC", x"FF", x"01", x"02", x"FF", x"FE", x"FE",
	x"FF", x"FE", x"FC", x"FC", x"FC", x"FB", x"F9", x"FB", x"FD", x"FD", x"FB", x"F9",
	x"F8", x"F9", x"FB", x"FB", x"FB", x"FA", x"F9", x"F9", x"FA", x"FB", x"FA", x"F8",
	x"F6", x"F7", x"F9", x"FC", x"FD", x"FD", x"FB", x"FB", x"FB", x"FA", x"FA", x"FC",
	x"FF", x"01", x"02", x"00", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FE", x"00", x"02", x"03",
	x"03", x"01", x"01", x"02", x"02", x"00", x"00", x"01", x"02", x"02", x"02", x"03",
	x"05", x"06", x"06", x"04", x"03", x"01", x"FF", x"00", x"02", x"04", x"03", x"02",
	x"03", x"03", x"02", x"01", x"02", x"04", x"04", x"02", x"03", x"03", x"03", x"03",
	x"03", x"02", x"01", x"01", x"01", x"02", x"03", x"04", x"03", x"FF", x"FC", x"FD",
	x"00", x"02", x"02", x"02", x"02", x"00", x"FE", x"FD", x"FE", x"FD", x"FC", x"FB",
	x"FB", x"FA", x"FB", x"FB", x"FC", x"FD", x"FD", x"FC", x"FA", x"FA", x"FA", x"FB",
	x"FD", x"FD", x"FD", x"FC", x"FB", x"FC", x"FB", x"F9", x"F8", x"FA", x"FD", x"00",
	x"00", x"FF", x"FC", x"FB", x"FC", x"FF", x"02", x"01", x"FF", x"FE", x"FF", x"00",
	x"02", x"02", x"01", x"00", x"01", x"01", x"00", x"00", x"01", x"04", x"04", x"02",
	x"01", x"01", x"02", x"04", x"04", x"05", x"05", x"05", x"06", x"05", x"03", x"03",
	x"02", x"01", x"01", x"01", x"03", x"04", x"03", x"01", x"FF", x"FD", x"FD", x"FF",
	x"00", x"00", x"00", x"01", x"02", x"01", x"FF", x"FE", x"FE", x"00", x"00", x"00",
	x"00", x"01", x"FF", x"FC", x"FA", x"F9", x"F8", x"F8", x"F9", x"F9", x"FA", x"FA",
	x"FA", x"FA", x"FC", x"FD", x"FC", x"FC", x"FD", x"FE", x"FE", x"FF", x"02", x"04",
	x"03", x"00", x"FE", x"FD", x"FD", x"FD", x"FE", x"00", x"02", x"03", x"03", x"01",
	x"FE", x"FC", x"FC", x"FE", x"01", x"01", x"00", x"00", x"01", x"02", x"01", x"01",
	x"01", x"01", x"00", x"FF", x"01", x"03", x"04", x"05", x"04", x"04", x"04", x"03",
	x"03", x"03", x"03", x"03", x"01", x"FF", x"FF", x"FE", x"FF", x"00", x"FE", x"FD",
	x"FD", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"FF", x"FD", x"FD", x"FE", x"FF",
	x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"FF",
	x"FD", x"FC", x"FC", x"FD", x"FD", x"FE", x"01", x"03", x"01", x"FF", x"FE", x"FE",
	x"FD", x"FA", x"F9", x"FB", x"FC", x"FB", x"FC", x"FD", x"FE", x"FD", x"FD", x"FD",
	x"FE", x"FC", x"FB", x"FA", x"FB", x"FB", x"FB", x"FC", x"FE", x"FD", x"FD", x"FC",
	x"FD", x"FD", x"FE", x"FF", x"FF", x"FE", x"FD", x"FD", x"FF", x"01", x"02", x"02",
	x"02", x"01", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"01", x"04", x"05", x"05",
	x"04", x"03", x"02", x"03", x"04", x"02", x"00", x"00", x"02", x"03", x"03", x"02",
	x"02", x"04", x"03", x"02", x"00", x"02", x"05", x"07", x"07", x"07", x"06", x"04",
	x"04", x"04", x"04", x"04", x"03", x"02", x"02", x"00", x"00", x"02", x"03", x"03",
	x"02", x"02", x"01", x"FF", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FD", x"FC", x"FB", x"FC", x"FC", x"FC", x"FD", x"FD", x"FC", x"FC", x"FD", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"FE", x"FD", x"FB", x"F8",
	x"F7", x"F7", x"FA", x"FC", x"FE", x"FD", x"FB", x"F9", x"F9", x"F9", x"F9", x"FA",
	x"FB", x"FC", x"FE", x"FF", x"FF", x"FF", x"01", x"01", x"00", x"FE", x"FE", x"FF",
	x"01", x"02", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"00",
	x"FE", x"FF", x"02", x"02", x"00", x"FE", x"FF", x"03", x"06", x"05", x"04", x"05",
	x"05", x"05", x"03", x"03", x"04", x"05", x"07", x"06", x"03", x"01", x"02", x"02",
	x"01", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FD", x"FE", x"FF", x"FE", x"FC",
	x"FB", x"FD", x"FE", x"FC", x"F9", x"F9", x"FC", x"FC", x"F9", x"F7", x"F9", x"FB",
	x"FB", x"FA", x"FA", x"FC", x"FD", x"FC", x"FA", x"F9", x"FA", x"FD", x"FE", x"FF",
	x"01", x"01", x"00", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE", x"FD", x"FE",
	x"00", x"00", x"FE", x"FF", x"03", x"05", x"03", x"02", x"02", x"03", x"04", x"04",
	x"03", x"03", x"05", x"05", x"05", x"06", x"07", x"07", x"05", x"03", x"03", x"04",
	x"04", x"05", x"05", x"05", x"05", x"04", x"04", x"04", x"03", x"03", x"02", x"02",
	x"01", x"02", x"03", x"02", x"FF", x"FE", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF",
	x"FE", x"FD", x"FD", x"FD", x"FB", x"F9", x"FA", x"FB", x"FC", x"FA", x"F9", x"FB",
	x"FC", x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FD", x"FC", x"FD", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE", x"FE", x"FF", x"00", x"02", x"05",
	x"05", x"02", x"FE", x"FD", x"FD", x"FE", x"FD", x"FD", x"FE", x"00", x"01", x"00",
	x"FE", x"FC", x"FC", x"FC", x"FB", x"FC", x"FD", x"FF", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FD", x"FC", x"FE", x"00", x"01", x"FE", x"FD", x"00", x"04", x"04", x"02",
	x"01", x"01", x"03", x"03", x"03", x"03", x"02", x"01", x"01", x"02", x"02", x"02",
	x"03", x"04", x"03", x"02", x"02", x"02", x"04", x"05", x"05", x"04", x"04", x"03",
	x"02", x"01", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"00", x"02", x"FF",
	x"FC", x"FB", x"FC", x"FC", x"FB", x"FA", x"FB", x"FA", x"FA", x"FA", x"FB", x"FE",
	x"FF", x"FD", x"FC", x"FA", x"FB", x"FE", x"FF", x"FE", x"FC", x"FE", x"00", x"FF",
	x"FE", x"FD", x"FD", x"FC", x"FA", x"F8", x"F9", x"FB", x"FC", x"FC", x"FD", x"FE",
	x"FD", x"FD", x"FE", x"00", x"01", x"02", x"02", x"00", x"FC", x"FA", x"FB", x"FE",
	x"00", x"FF", x"FD", x"FE", x"00", x"00", x"FF", x"FF", x"FD", x"FC", x"FC", x"FD",
	x"FF", x"00", x"01", x"03", x"04", x"03", x"01", x"FE", x"FD", x"FD", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"01", x"03", x"02", x"00", x"01", x"05", x"06",
	x"05", x"04", x"05", x"06", x"06", x"06", x"06", x"08", x"0A", x"08", x"05", x"03",
	x"02", x"01", x"02", x"02", x"03", x"02", x"00", x"FD", x"FC", x"FC", x"FD", x"FC",
	x"FA", x"FB", x"FC", x"FC", x"FB", x"FC", x"FE", x"00", x"FF", x"FC", x"FB", x"FC",
	x"FE", x"FE", x"FE", x"01", x"02", x"FF", x"FE", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FD", x"FC", x"FD", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FD", x"FC",
	x"FD", x"00", x"02", x"00", x"FF", x"00", x"02", x"03", x"03", x"03", x"03", x"03",
	x"04", x"04", x"04", x"03", x"02", x"02", x"02", x"03", x"04", x"06", x"07", x"07",
	x"06", x"05", x"04", x"02", x"01", x"01", x"03", x"03", x"01", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"01", x"02", x"03", x"02", x"00", x"FD", x"FC", x"FC", x"FA",
	x"F8", x"F8", x"FA", x"FB", x"FA", x"FA", x"FA", x"FB", x"FC", x"FB", x"FB", x"FA",
	x"FA", x"FA", x"FA", x"FC", x"FE", x"FE", x"FC", x"FB", x"FA", x"F9", x"F9", x"FB",
	x"FD", x"FB", x"FB", x"FC", x"FC", x"FC", x"FA", x"FB", x"FD", x"FC", x"FC", x"FC",
	x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"FF", x"FE", x"FF", x"00",
	x"00", x"01", x"01", x"00", x"01", x"02", x"03", x"04", x"03", x"01", x"00", x"00",
	x"01", x"01", x"FF", x"00", x"00", x"00", x"FF", x"01", x"03", x"03", x"02", x"01",
	x"FF", x"FF", x"FF", x"00", x"01", x"01", x"FF", x"FD", x"FE", x"01", x"02", x"00",
	x"00", x"02", x"04", x"05", x"04", x"03", x"03", x"03", x"03", x"03", x"03", x"03",
	x"02", x"01", x"00", x"00", x"01", x"01", x"01", x"02", x"03", x"01", x"00", x"00",
	x"02", x"02", x"02", x"01", x"01", x"FF", x"FE", x"FD", x"FE", x"00", x"00", x"FF",
	x"FE", x"FD", x"FC", x"FB", x"FB", x"FA", x"FA", x"F9", x"F9", x"FE", x"03", x"03",
	x"02", x"00", x"00", x"00", x"FF", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FC", x"FA", x"FA", x"F8", x"F8", x"FB", x"FF", x"FE", x"FA", x"FA", x"FD",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"04", x"05", x"06", x"05", x"04", x"03", x"01", x"01", x"02",
	x"02", x"02", x"01", x"00", x"FF", x"00", x"00", x"01", x"01", x"03", x"05", x"04",
	x"03", x"01", x"00", x"01", x"01", x"FF", x"FF", x"01", x"03", x"04", x"03", x"01",
	x"01", x"01", x"01", x"FF", x"FE", x"FE", x"FE", x"FE", x"FD", x"FB", x"FA", x"FB",
	x"FC", x"FB", x"FA", x"FB", x"FC", x"FB", x"FB", x"FA", x"FB", x"FC", x"FC", x"FD",
	x"FE", x"00", x"FF", x"FD", x"FD", x"FD", x"FC", x"FB", x"FC", x"FD", x"FD", x"FD",
	x"FD", x"FE", x"FF", x"FF", x"FF", x"01", x"02", x"00", x"FE", x"FE", x"FE", x"FE",
	x"FD", x"FE", x"FF", x"FE", x"FC", x"FC", x"FF", x"00", x"FF", x"FF", x"00", x"00",
	x"FF", x"01", x"03", x"04", x"03", x"02", x"03", x"05", x"06", x"04", x"03", x"04",
	x"06", x"06", x"05", x"04", x"05", x"06", x"05", x"05", x"06", x"06", x"05", x"03",
	x"03", x"03", x"03", x"03", x"03", x"02", x"01", x"00", x"00", x"00", x"00", x"00",
	x"FE", x"FD", x"FC", x"FD", x"FC", x"FC", x"FE", x"FF", x"FE", x"FB", x"F9", x"F8",
	x"FA", x"FD", x"FD", x"FC", x"FB", x"FB", x"FA", x"F9", x"FA", x"FA", x"F8", x"F8",
	x"F9", x"F8", x"F5", x"F6", x"F9", x"FA", x"FC", x"FC", x"FC", x"FB", x"FB", x"FC",
	x"FD", x"FE", x"00", x"00", x"FF", x"FE", x"FD", x"FD", x"FF", x"02", x"03", x"00",
	x"FE", x"FE", x"00", x"01", x"FF", x"FF", x"02", x"05", x"05", x"04", x"05", x"07",
	x"07", x"06", x"07", x"06", x"04", x"02", x"03", x"04", x"04", x"05", x"07", x"08",
	x"05", x"02", x"02", x"02", x"02", x"02", x"03", x"04", x"03", x"02", x"01", x"00",
	x"00", x"00", x"01", x"02", x"02", x"02", x"01", x"01", x"01", x"00", x"FF", x"FE",
	x"FD", x"FD", x"00", x"01", x"01", x"FF", x"FD", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FD", x"FE", x"FE", x"FD", x"FE", x"FF", x"FF", x"FE", x"FD", x"FC", x"FC", x"FE",
	x"FF", x"FF", x"FE", x"FD", x"FD", x"FE", x"FE", x"FD", x"FC", x"FC", x"FD", x"FD",
	x"FD", x"FD", x"FE", x"00", x"01", x"00", x"FF", x"FE", x"00", x"01", x"00", x"00",
	x"01", x"00", x"FF", x"FC", x"FA", x"FA", x"FD", x"FE", x"FC", x"FA", x"FA", x"FA",
	x"F9", x"F7", x"F7", x"FA", x"FB", x"FB", x"FB", x"FB", x"FE", x"00", x"01", x"01",
	x"02", x"03", x"04", x"04", x"04", x"04", x"05", x"06", x"04", x"03", x"03", x"03",
	x"03", x"03", x"02", x"01", x"01", x"01", x"01", x"02", x"03", x"03", x"02", x"01",
	x"00", x"01", x"03", x"04", x"03", x"02", x"01", x"01", x"01", x"01", x"00", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FC", x"FB", x"FB", x"FC",
	x"FC", x"FB", x"FB", x"FC", x"FD", x"FD", x"FD", x"FD", x"FF", x"FE", x"FD", x"FC",
	x"FC", x"FD", x"FC", x"FB", x"FA", x"FC", x"FC", x"FC", x"FD", x"FE", x"FF", x"00",
	x"FF", x"FE", x"FF", x"01", x"01", x"00", x"FF", x"FE", x"00", x"03", x"03", x"00",
	x"FF", x"00", x"FF", x"FE", x"FD", x"FE", x"00", x"00", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"01", x"03", x"03", x"02", x"03", x"05", x"06", x"06", x"05", x"04",
	x"03", x"02", x"03", x"04", x"04", x"03", x"02", x"01", x"02", x"03", x"02", x"02",
	x"02", x"02", x"03", x"02", x"01", x"00", x"01", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FD", x"FE", x"00", x"00", x"FF", x"FD", x"FD", x"FC", x"FB", x"F9",
	x"F8", x"F8", x"F8", x"F9", x"FB", x"FD", x"FD", x"FC", x"FC", x"FE", x"FE", x"FE",
	x"FD", x"FD", x"FE", x"FE", x"FD", x"FC", x"FD", x"FE", x"FE", x"FD", x"FD", x"FE",
	x"FD", x"FD", x"FD", x"FD", x"FC", x"FA", x"FB", x"FC", x"FC", x"FB", x"FD", x"FF",
	x"02", x"03", x"03", x"03", x"03", x"02", x"00", x"FF", x"FF", x"FF", x"00", x"02",
	x"05", x"07", x"06", x"04", x"04", x"05", x"05", x"04", x"02", x"02", x"02", x"01",
	x"02", x"05", x"06", x"06", x"03", x"02", x"03", x"03", x"02", x"02", x"02", x"02",
	x"02", x"02", x"01", x"00", x"FF", x"FE", x"FE", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FD", x"FD", x"FE", x"FD", x"FC", x"FC", x"FD", x"FE", x"FD", x"FD",
	x"FD", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FC", x"FB", x"FB", x"FD", x"FE",
	x"FD", x"FD", x"FE", x"FF", x"FE", x"FE", x"00", x"00", x"FD", x"FD", x"FE", x"FF",
	x"00", x"00", x"00", x"01", x"02", x"03", x"02", x"00", x"00", x"00", x"01", x"02",
	x"FF", x"FE", x"FE", x"FE", x"FC", x"FA", x"FB", x"FC", x"FD", x"FE", x"FD", x"FD",
	x"FD", x"FE", x"FD", x"FC", x"FD", x"FE", x"FD", x"FB", x"FA", x"FA", x"FA", x"FB",
	x"FB", x"FD", x"FF", x"00", x"00", x"FF", x"00", x"01", x"01", x"02", x"02", x"03",
	x"02", x"00", x"FF", x"00", x"02", x"03", x"04", x"07", x"07", x"05", x"03", x"03",
	x"02", x"02", x"01", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF",
	x"00", x"01", x"02", x"02", x"01", x"01", x"00", x"01", x"01", x"02", x"01", x"00",
	x"FF", x"FF", x"FF", x"FD", x"FC", x"FC", x"FC", x"FC", x"FD", x"FD", x"FD", x"FC",
	x"FB", x"FA", x"FA", x"F9", x"F9", x"FA", x"FC", x"FC", x"FA", x"FA", x"FB", x"FE",
	x"00", x"FF", x"FC", x"FB", x"FB", x"FC", x"FB", x"FD", x"FF", x"FF", x"FD", x"FE",
	x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"03", x"03", x"02", x"01",
	x"01", x"00", x"00", x"01", x"03", x"04", x"04", x"04", x"03", x"04", x"04", x"04",
	x"03", x"03", x"04", x"05", x"05", x"04", x"03", x"05", x"06", x"05", x"03", x"02",
	x"01", x"01", x"01", x"00", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FE", x"FD", x"FE", x"FF", x"FE", x"FC", x"FA", x"F8", x"F8", x"FA",
	x"FB", x"FC", x"FC", x"FD", x"FC", x"FB", x"FA", x"FB", x"FD", x"FE", x"FE", x"FD",
	x"FD", x"FE", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FC", x"FD", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FD", x"FC", x"FD", x"FE", x"FE", x"FD", x"FD", x"FF",
	x"00", x"00", x"00", x"01", x"00", x"FE", x"FE", x"00", x"01", x"01", x"00", x"00",
	x"01", x"02", x"03", x"03", x"03", x"04", x"05", x"06", x"06", x"04", x"02", x"02",
	x"02", x"02", x"03", x"03", x"02", x"03", x"05", x"04", x"01", x"00", x"01", x"01",
	x"01", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FE", x"FD", x"FC", x"FD", x"FE", x"FE", x"FD", x"FD", x"FE", x"FE",
	x"FE", x"FE", x"FD", x"FB", x"FB", x"FD", x"FD", x"FC", x"FC", x"FE", x"FE", x"FC",
	x"FB", x"FB", x"FC", x"FD", x"FF", x"01", x"01", x"00", x"FF", x"FE", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"03", x"04", x"04", x"03",
	x"01", x"01", x"02", x"01", x"01", x"01", x"01", x"00", x"00", x"01", x"01", x"00",
	x"FF", x"FF", x"00", x"01", x"FF", x"FD", x"FD", x"FE", x"FF", x"FE", x"FD", x"FF",
	x"01", x"02", x"01", x"01", x"02", x"02", x"03", x"02", x"02", x"01", x"01", x"00",
	x"00", x"03", x"03", x"03", x"03", x"02", x"00", x"FE", x"FD", x"FF", x"00", x"00",
	x"00", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FE", x"FD", x"FC", x"FB", x"FC", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FF", x"00", x"00", x"FE", x"FB", x"FA", x"F9", x"F9", x"F9", x"FA", x"FA", x"F9",
	x"F8", x"F8", x"F8", x"F9", x"FA", x"FA", x"FC", x"FE", x"00", x"00", x"02", x"03",
	x"01", x"FE", x"FD", x"FE", x"00", x"01", x"02", x"04", x"04", x"02", x"01", x"01",
	x"01", x"00", x"FF", x"00", x"02", x"03", x"04", x"03", x"03", x"04", x"05", x"05",
	x"03", x"02", x"03", x"03", x"03", x"02", x"05", x"07", x"06", x"04", x"03", x"03",
	x"02", x"00", x"FF", x"FF", x"FD", x"FA", x"F9", x"FA", x"FB", x"FC", x"FD", x"FF",
	x"FF", x"FD", x"FC", x"FC", x"FC", x"FB", x"FA", x"FA", x"FB", x"FD", x"FE", x"FE",
	x"FD", x"FD", x"FE", x"FE", x"FD", x"FC", x"FD", x"FC", x"FB", x"FB", x"FB", x"FB",
	x"FC", x"FE", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"03", x"02", x"01",
	x"00", x"01", x"01", x"01", x"01", x"02", x"03", x"03", x"02", x"01", x"00", x"00",
	x"00", x"00", x"00", x"01", x"01", x"02", x"03", x"03", x"01", x"01", x"02", x"03",
	x"02", x"03", x"05", x"04", x"03", x"02", x"01", x"01", x"01", x"01", x"02", x"02",
	x"02", x"03", x"03", x"03", x"03", x"02", x"01", x"02", x"03", x"01", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FD",
	x"FC", x"FB", x"FA", x"FA", x"FC", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"00",
	x"FF", x"FD", x"FC", x"FC", x"FD", x"FE", x"FE", x"FE", x"FE", x"FF", x"FE", x"FC",
	x"FC", x"FD", x"FE", x"FD", x"FC", x"FB", x"FC", x"FD", x"FC", x"FD", x"FE", x"00",
	x"01", x"00", x"01", x"02", x"01", x"FF", x"FE", x"FF", x"00", x"FF", x"FE", x"FE",
	x"01", x"04", x"04", x"02", x"01", x"01", x"01", x"00", x"FF", x"00", x"01", x"01",
	x"00", x"FE", x"FF", x"FF", x"FF", x"01", x"02", x"02", x"01", x"01", x"02", x"02",
	x"02", x"02", x"02", x"02", x"01", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FC", x"FD", x"FE", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FF", x"FF", x"FE", x"FD", x"FD",
	x"FC", x"FB", x"FA", x"FA", x"FA", x"FB", x"FC", x"FD", x"FD", x"FC", x"FB", x"FD",
	x"FF", x"00", x"01", x"04", x"03", x"00", x"FC", x"FB", x"FD", x"FF", x"00", x"01",
	x"02", x"01", x"FF", x"FE", x"FF", x"FE", x"FC", x"FA", x"FA", x"FB", x"FB", x"FC",
	x"FD", x"FE", x"FF", x"00", x"00", x"FF", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"01", x"00",
	x"00", x"02", x"03", x"03", x"02", x"02", x"02", x"02", x"03", x"03", x"04", x"04",
	x"03", x"03", x"03", x"04", x"03", x"03", x"05", x"06", x"06", x"05", x"06", x"07",
	x"06", x"05", x"05", x"04", x"03", x"02", x"03", x"02", x"02", x"01", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"FF", x"FD", x"FD", x"FE", x"FD",
	x"FD", x"FE", x"FE", x"FD", x"FA", x"F8", x"FA", x"FB", x"FA", x"FA", x"FB", x"FD",
	x"FC", x"F9", x"F7", x"F8", x"FA", x"F9", x"FB", x"FE", x"01", x"01", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"01",
	x"02", x"02", x"00", x"FF", x"FF", x"01", x"01", x"01", x"03", x"03", x"02", x"01",
	x"01", x"02", x"01", x"01", x"02", x"03", x"03", x"01", x"FF", x"00", x"02", x"02",
	x"02", x"01", x"00", x"FE", x"FC", x"FC", x"FE", x"00", x"02", x"03", x"02", x"01",
	x"00", x"00", x"FF", x"FD", x"FC", x"FC", x"FC", x"FC", x"FD", x"FF", x"00", x"FF",
	x"FF", x"FE", x"FD", x"FE", x"FE", x"FD", x"FD", x"FD", x"FC", x"FC", x"FD", x"FE",
	x"FE", x"FD", x"FC", x"FC", x"FD", x"FD", x"FD", x"FC", x"FB", x"FC", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FE", x"FF", x"FE", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FE", x"FF", x"00", x"01", x"01", x"00", x"00", x"01", x"01", x"00",
	x"00", x"00", x"FF", x"FE", x"FF", x"02", x"04", x"03", x"01", x"00", x"FE", x"FF",
	x"00", x"01", x"01", x"01", x"01", x"02", x"04", x"04", x"05", x"05", x"04", x"04",
	x"05", x"06", x"05", x"04", x"03", x"03", x"02", x"00", x"FF", x"00", x"00", x"00",
	x"01", x"01", x"02", x"02", x"02", x"01", x"01", x"02", x"02", x"02", x"02", x"03",
	x"02", x"01", x"00", x"00", x"00", x"FF", x"FD", x"FC", x"FC", x"FC", x"FD", x"FF",
	x"FE", x"FD", x"FB", x"FC", x"FE", x"FE", x"FD", x"FD", x"FE", x"FD", x"FB", x"FB",
	x"FC", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE",
	x"FC", x"FE", x"00", x"01", x"01", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"01",
	x"02", x"01", x"FF", x"FE", x"FE", x"FF", x"01", x"01", x"00", x"01", x"02", x"01",
	x"00", x"FF", x"00", x"01", x"01", x"00", x"FF", x"FF", x"00", x"01", x"00", x"00",
	x"00", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"00", x"01", x"00", x"FF", x"FD", x"FD", x"FE", x"FD", x"FE", x"00", x"01",
	x"01", x"00", x"FF", x"FF", x"FE", x"FD", x"FC", x"FB", x"FA", x"F9", x"F9", x"FB",
	x"FE", x"FF", x"00", x"FF", x"FD", x"FC", x"FC", x"FC", x"FB", x"FC", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"FE", x"FC", x"FC", x"FE", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"02", x"01", x"01", x"FF",
	x"FE", x"FE", x"00", x"01", x"02", x"03", x"03", x"03", x"02", x"03", x"03", x"02",
	x"01", x"02", x"02", x"02", x"01", x"02", x"04", x"04", x"03", x"01", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FD", x"FB", x"FB", x"FB", x"FB", x"FC",
	x"FD", x"FE", x"FE", x"FD", x"FD", x"FE", x"FE", x"FD", x"FD", x"FE", x"FE", x"FD",
	x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"02", x"01", x"00", x"FF",
	x"FE", x"FD", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"00", x"01", x"00", x"FE",
	x"FE", x"FF", x"FF", x"00", x"02", x"03", x"04", x"04", x"04", x"04", x"03", x"02",
	x"00", x"00", x"FF", x"00", x"01", x"02", x"02", x"02", x"02", x"02", x"02", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"02", x"02", x"02", x"01", x"01", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FE", x"FE", x"00", x"02", x"01",
	x"FF", x"FE", x"FD", x"FC", x"FD", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FE", x"FC", x"FB", x"FC", x"FD", x"FE", x"FE", x"FF", x"FF",
	x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FB", x"FB", x"FC", x"FE", x"FE", x"FD",
	x"FD", x"FD", x"FD", x"FC", x"FC", x"FD", x"FD", x"FD", x"FE", x"FF", x"00", x"FE",
	x"FC", x"FB", x"FE", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"01", x"02", x"02", x"02", x"02", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01",
	x"02", x"02", x"02", x"01", x"00", x"FF", x"00", x"01", x"03", x"04", x"04", x"03",
	x"03", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01",
	x"00", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FD", x"FE",
	x"00", x"03", x"03", x"01", x"00", x"FF", x"FE", x"FD", x"FD", x"FE", x"00", x"01",
	x"01", x"01", x"01", x"00", x"00", x"01", x"03", x"03", x"02", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FE", x"FC", x"FD",
	x"FE", x"FD", x"FD", x"FD", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE",
	x"FE", x"FE", x"FD", x"FE", x"FF", x"FE", x"FD", x"FD", x"FE", x"FF", x"01", x"02",
	x"01", x"00", x"00", x"02", x"01", x"01", x"02", x"04", x"04", x"03", x"01", x"00",
	x"FF", x"00", x"FF", x"00", x"01", x"02", x"02", x"01", x"FF", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FE", x"FE", x"FD", x"FB", x"FB", x"FD", x"FD", x"FD", x"FD", x"FE",
	x"FF", x"FD", x"FC", x"FC", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FB", x"FA",
	x"FC", x"FF", x"FE", x"FD", x"FE", x"FF", x"FE", x"FD", x"FC", x"FD", x"FE", x"FE",
	x"FE", x"FE", x"00", x"00", x"01", x"01", x"01", x"02", x"02", x"02", x"02", x"02",
	x"01", x"01", x"01", x"02", x"01", x"02", x"03", x"04", x"04", x"03", x"03", x"04",
	x"05", x"04", x"03", x"02", x"01", x"00", x"FF", x"00", x"02", x"02", x"02", x"01",
	x"01", x"00", x"FF", x"FF", x"FF", x"01", x"02", x"02", x"01", x"00", x"00", x"02",
	x"02", x"01", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FC", x"FC", x"FC",
	x"FC", x"FC", x"FD", x"FD", x"FE", x"FE", x"FD", x"FC", x"FC", x"FC", x"FD", x"FD",
	x"FE", x"FF", x"FF", x"FE", x"FD", x"FD", x"FC", x"FB", x"FB", x"FD", x"FE", x"FE",
	x"FE", x"FF", x"01", x"01", x"01", x"00", x"FF", x"FF", x"00", x"01", x"00", x"FF",
	x"FF", x"FF", x"00", x"01", x"02", x"02", x"02", x"01", x"01", x"01", x"00", x"FF",
	x"FF", x"01", x"01", x"FF", x"FF", x"00", x"FE", x"FC", x"FC", x"FF", x"01", x"02",
	x"03", x"03", x"02", x"02", x"02", x"03", x"03", x"02", x"02", x"02", x"03", x"02",
	x"01", x"01", x"03", x"03", x"01", x"FF", x"FF", x"FF", x"FF", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FC", x"FD", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FE",
	x"FF", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FD",
	x"FC", x"FD", x"FE", x"FF", x"FF", x"00", x"01", x"00", x"00", x"01", x"02", x"02",
	x"02", x"00", x"FF", x"FE", x"FE", x"FD", x"FC", x"FD", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FD", x"FD", x"FD", x"FE", x"00",
	x"01", x"02", x"02", x"02", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FE", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FD",
	x"FE", x"FF", x"FF", x"FE", x"FF", x"02", x"03", x"03", x"02", x"01", x"01", x"02",
	x"01", x"01", x"01", x"02", x"02", x"02", x"02", x"01", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FE", x"FD", x"FD", x"FD",
	x"FD", x"FC", x"FC", x"FC", x"FB", x"FB", x"FC", x"FC", x"FC", x"FC", x"FD", x"FE",
	x"FE", x"FD", x"FC", x"FC", x"FD", x"FE", x"FE", x"FE", x"FF", x"00", x"FF", x"FE",
	x"FF", x"00", x"01", x"01", x"02", x"02", x"01", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"01", x"02", x"03", x"04", x"03", x"02", x"01", x"01", x"01", x"02",
	x"03", x"04", x"04", x"04", x"03", x"02", x"03", x"04", x"04", x"03", x"02", x"01",
	x"FF", x"FE", x"FF", x"00", x"00", x"01", x"00", x"01", x"01", x"01", x"01", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FD", x"FB", x"FA", x"F9", x"F9", x"FA", x"FB", x"FB", x"FB", x"FB", x"FC", x"FC",
	x"FC", x"FD", x"FD", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FE", x"FD", x"FD",
	x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"00", x"00",
	x"00", x"FF", x"FE", x"FF", x"00", x"02", x"01", x"01", x"01", x"02", x"02", x"02",
	x"02", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"02", x"03",
	x"03", x"02", x"02", x"03", x"03", x"01", x"00", x"01", x"01", x"00", x"00", x"00",
	x"01", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FE", x"FE", x"00", x"02",
	x"02", x"01", x"01", x"01", x"FF", x"FE", x"FD", x"FE", x"FF", x"FF", x"FE", x"FF",
	x"00", x"01", x"00", x"00", x"00", x"FF", x"FD", x"FD", x"FF", x"01", x"01", x"01",
	x"02", x"01", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FD", x"FD", x"FE", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FD", x"FD", x"FD", x"FF",
	x"FF", x"FF", x"FE", x"FD", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"01", x"03", x"04", x"04",
	x"02", x"00", x"00", x"01", x"02", x"02", x"01", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"02", x"02", x"01", x"FF", x"FD", x"FC", x"FC", x"FC", x"FD", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FD", x"FD", x"FD", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF",
	x"FE", x"FD", x"FD", x"FE", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"01", x"01", x"00", x"00",
	x"02", x"02", x"01", x"01", x"02", x"02", x"02", x"02", x"04", x"05", x"04", x"03",
	x"03", x"03", x"02", x"02", x"03", x"03", x"02", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"01", x"02", x"02", x"01", x"00", x"00", x"00", x"FE",
	x"FD", x"FC", x"FC", x"FD", x"FD", x"FC", x"FB", x"FB", x"FC", x"FC", x"FA", x"FA",
	x"FC", x"FC", x"FA", x"F9", x"F9", x"FA", x"FB", x"FB", x"FC", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"00", x"01",
	x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"02", x"02", x"02", x"02", x"01", x"02", x"02", x"01", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"01", x"00", x"FF", x"FE", x"FD", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"00", x"01",
	x"02", x"02", x"02", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02",
	x"03", x"02", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"01", x"01", x"01", x"01", x"00",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"00", x"02", x"03", x"02", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"00", x"FF", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FE", x"FE", x"FF", x"00",
	x"00", x"01", x"02", x"03", x"02", x"01", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"02",
	x"02", x"01", x"FF", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"00", x"02", x"01", x"FF", x"FF", x"00", x"FF", x"FE", x"FD", x"FE", x"FE", x"FF",
	x"FF", x"00", x"01", x"02", x"01", x"00", x"00", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"01", x"00", x"FF", x"FE", x"FF", x"00", x"01", x"01", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"00",
	x"01", x"01", x"00", x"00", x"01", x"02", x"01", x"01", x"00", x"00", x"00", x"01",
	x"01", x"01", x"01", x"01", x"01", x"00", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE", x"FE", x"FE", x"FD",
	x"FD", x"FC", x"FC", x"FB", x"FA", x"F9", x"FA", x"FB", x"FD", x"FD", x"FC", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"02", x"02", x"02", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"01", x"00", x"FF", x"FF", x"01", x"02", x"02", x"01", x"00", x"FF", x"FF", x"00",
	x"00", x"02", x"02", x"02", x"01", x"00", x"01", x"01", x"02", x"02", x"01", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FE", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FE", x"FD",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"00", x"FF", x"FE", x"FE", x"FF", x"01", x"02", x"02", x"02", x"01", x"FF", x"FE",
	x"FE", x"FF", x"FF", x"00", x"01", x"02", x"03", x"02", x"02", x"02", x"01", x"FF",
	x"FF", x"01", x"02", x"03", x"03", x"02", x"01", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FD", x"FC", x"FC", x"FC", x"FD", x"FC", x"FB", x"FC", x"FE", x"FF",
	x"FF", x"FE", x"FE", x"FC", x"FB", x"FB", x"FC", x"FE", x"FF", x"00", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"00", x"00", x"FF",
	x"00", x"01", x"00", x"FF", x"FE", x"FF", x"00", x"FE", x"FE", x"FF", x"00", x"01",
	x"00", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"00", x"01", x"01",
	x"01", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FD",
	x"FD", x"FD", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FD",
	x"FC", x"FC", x"FD", x"FE", x"FE", x"FD", x"FD", x"FE", x"FF", x"00", x"00", x"01",
	x"01", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"01", x"01", x"00", x"00",
	x"01", x"02", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"02",
	x"02", x"01", x"00", x"FF", x"FF", x"00", x"01", x"02", x"01", x"01", x"01", x"02",
	x"02", x"02", x"01", x"01", x"01", x"01", x"02", x"01", x"01", x"00", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"FD", x"FC", x"FD", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FC", x"FC", x"FD", x"FD",
	x"FD", x"FE", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"FF",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FD", x"FC",
	x"FD", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"02", x"04", x"04", x"03",
	x"03", x"03", x"02", x"01", x"01", x"01", x"02", x"02", x"02", x"01", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"00", x"FF", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE", x"FE", x"FD", x"FC", x"FC",
	x"FC", x"FC", x"FC", x"FC", x"FD", x"FD", x"FD", x"FE", x"FF", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"03", x"03",
	x"03", x"01", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"FE", x"FE", x"FE", x"FD",
	x"FC", x"FC", x"FC", x"FE", x"FE", x"FD", x"FD", x"FE", x"00", x"01", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"01", x"01", x"01",
	x"02", x"02", x"02", x"02", x"02", x"03", x"03", x"02", x"02", x"03", x"03", x"02",
	x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"01",
	x"01", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FC", x"FD", x"FE", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"02", x"01", x"01", x"02",
	x"03", x"03", x"03", x"03", x"03", x"01", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FE", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00",
	x"01", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"01", x"02", x"02",
	x"01", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD",
	x"FC", x"FC", x"FD", x"FD", x"FC", x"FC", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE",
	x"FD", x"FD", x"FD", x"FD", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"01", x"02", x"01",
	x"00", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"00",
	x"01", x"02", x"02", x"02", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01",
	x"00", x"00", x"01", x"02", x"02", x"01", x"01", x"02", x"02", x"01", x"00", x"00",
	x"01", x"02", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FD", x"FE", x"FE", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD",
	x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"FD",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00",
	x"02", x"03", x"02", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"00", x"00",
	x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"01", x"00", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"02", x"02", x"02", x"01", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01",
	x"00", x"00", x"00", x"01", x"02", x"01", x"00", x"FF", x"FE", x"FE", x"FD", x"FD",
	x"FE", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FE",
	x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE",
	x"FE", x"FC", x"FB", x"FC", x"FD", x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"01",
	x"01", x"02", x"03", x"04", x"04", x"03", x"03", x"02", x"03", x"03", x"03", x"03",
	x"03", x"01", x"00", x"00", x"00", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"02", x"02", x"02", x"01", x"FE",
	x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"02", x"03", x"03", x"02", x"02", x"01",
	x"01", x"00", x"00", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD",
	x"FE", x"00", x"00", x"01", x"01", x"00", x"01", x"02", x"02", x"02", x"02", x"02",
	x"02", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FE", x"FD", x"FD", x"FE", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FE", x"FD", x"FC", x"FB", x"FB", x"FC", x"FD", x"FD", x"FE", x"FE",
	x"FE", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"01", x"01", x"00", x"00", x"00", x"01", x"00", x"FF", x"FF", x"00", x"00",
	x"FF", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"00",
	x"02", x"02", x"01", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"02", x"01", x"00", x"FF", x"FF", x"00", x"00", x"FF",
	x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FC", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"01", x"01", x"01", x"02", x"02", x"01", x"01", x"01", x"02",
	x"01", x"01", x"02", x"02", x"02", x"02", x"02", x"02", x"00", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FD", x"FC", x"FD", x"FE", x"FE", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FD", x"FC", x"FD", x"FE", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"02", x"02", x"01", x"FF",
	x"FE", x"FE", x"FF", x"00", x"00", x"00", x"01", x"02", x"02", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"01", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FD",
	x"FD", x"FE", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FD", x"FD", x"FF", x"00",
	x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE",
	x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"01", x"00", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF",
	x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FC",
	x"FD", x"FE", x"FE", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FE", x"FE",
	x"FF", x"00", x"00", x"FF", x"00", x"01", x"01", x"01", x"00", x"01", x"01", x"01",
	x"01", x"00", x"00", x"00", x"01", x"00", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"02", x"02", x"01", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"00", x"00", x"FF", x"FF", x"00", x"01", x"02", x"03", x"02", x"01", x"01", x"00",
	x"FF", x"FF", x"01", x"02", x"02", x"02", x"02", x"02", x"01", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"FF", x"FE", x"FD", x"FC", x"FD", x"FE", x"FE", x"FD",
	x"FD", x"FD", x"FD", x"FB", x"FA", x"FB", x"FC", x"FD", x"FC", x"FB", x"FB", x"FD",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"01", x"02", x"01", x"01", x"01", x"01", x"00",
	x"00", x"FF", x"00", x"00", x"01", x"00", x"00", x"01", x"02", x"03", x"03", x"02",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FE", x"FD", x"FD", x"FE",
	x"FF", x"FF", x"FD", x"FC", x"FD", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00",
	x"01", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"00", x"00", x"FF", x"FE", x"FE", x"FD", x"FE", x"FF", x"01", x"01", x"01",
	x"00", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FD",
	x"FD", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00",
	x"FF", x"FE", x"FD", x"FD", x"FD", x"FF", x"00", x"01", x"FF", x"FE", x"FE", x"FE",
	x"FD", x"FD", x"FC", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"01", x"01", x"02", x"02", x"03",
	x"03", x"03", x"03", x"03", x"01", x"00", x"00", x"00", x"01", x"02", x"01", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE", x"FE", x"FD", x"FE", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"FD", x"FC", x"FC", x"FD",
	x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FE", x"FF", x"00", x"01", x"03", x"03", x"02", x"01",
	x"01", x"02", x"03", x"03", x"02", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00",
	x"01", x"01", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FD", x"FC", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FE", x"FF", x"FF", x"FE", x"FD", x"FD", x"FE", x"FE", x"FD", x"FD", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"00", x"01",
	x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"00", x"01", x"02", x"01", x"00",
	x"01", x"01", x"02", x"03", x"03", x"02", x"01", x"00", x"00", x"01", x"01", x"00",
	x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"01", x"01", x"01", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FE",
	x"FD", x"FD", x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"FF", x"FE", x"FE", x"FD",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FD", x"FE", x"FF", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"01", x"00", x"01",
	x"01", x"00", x"00", x"01", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"01", x"02", x"02", x"02", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FC", x"FD", x"FE", x"FF", x"00",
	x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"01", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FE", x"FD", x"FD",
	x"FE", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FD", x"FC", x"FC",
	x"FD", x"FD", x"FC", x"FC", x"FC", x"FD", x"FD", x"FC", x"FC", x"FD", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"01", x"01", x"01", x"01", x"03", x"03", x"02", x"02",
	x"01", x"00", x"01", x"01", x"01", x"00", x"01", x"02", x"01", x"01", x"00", x"01",
	x"00", x"00", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"01",
	x"01", x"01", x"02", x"02", x"00", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FE",
	x"FE", x"FD", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00",
	x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"02", x"02", x"02", x"02",
	x"02", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"02", x"02", x"01", x"01",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"00", x"01",
	x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"01", x"02", x"02", x"02", x"02", x"01", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"01", x"01", x"01", x"00", x"00", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"02", x"02", x"01", x"01", x"01",
	x"00", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"02", x"02", x"03", x"02", x"02",
	x"02", x"02", x"02", x"02", x"01", x"00", x"00", x"01", x"01", x"02", x"02", x"02",
	x"01", x"01", x"01", x"01", x"00", x"FF", x"00", x"00", x"FF", x"FE", x"FD", x"FD",
	x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD",
	x"FD", x"FC", x"FC", x"FD", x"FD", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"02", x"02", x"01", x"01",
	x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"01", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"01", x"01", x"00", x"FF", x"00", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FD", x"FD",
	x"FE", x"FF", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"00", x"01", x"01", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"01", x"01",
	x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00",
	x"01", x"01", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FD", x"FD", x"FE", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"01", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"01", x"01",
	x"01", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"01", x"01", x"02", x"01", x"01", x"01", x"01", x"01", x"00",
	x"01", x"02", x"02", x"02", x"02", x"01", x"00", x"00", x"00", x"00", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FC", x"FC", x"FD", x"FD", x"FE",
	x"FE"
	);

	
signal cnt_out: integer := 0;	
signal play_sound: std_logic := '0';
constant cnt_max: integer := 19213;
--signal out_signal: signed(7 downto 0) := x"00";

begin
	
process (CLK)
begin
    if rising_edge(CLK) then
        if RST = '1' then
            play_sound <= '0';
        elsif PLAY = '1' then
            play_sound <= '1';
        elsif PLAY = '0' and cnt_out = cnt_max then
            play_sound <= '0';
        end if;
    end if;
end process;

	
--counter
process (CLK)
begin     
    if rising_edge(CLK) then
        if RST = '1' then
            cnt_out <= 0;
        elsif CE = '1' and play_sound = '1' then
            cnt_out <= cnt_out + 1;       
        end if;
        if cnt_out = cnt_max then
            cnt_out <= 0;            
        end if;        
    end if;
end process;

process (CLK) 
begin
    if rising_edge(CLK) then
        if RST = '1' then
            SNARE_SAMP_O <= x"00";
        elsif CE = '1' then
            SNARE_SAMP_O <= snare_sound(cnt_out);
        end if;
    end if;    
end process;

end Behavioral;