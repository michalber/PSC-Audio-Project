----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 25.12.2018 17:39:59
-- Design Name: 
-- Module Name: Tom2 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Tom2 is
    Port ( CLK : in STD_LOGIC;
           CE : in STD_LOGIC;
           RST : in STD_LOGIC;
           PLAY : in STD_LOGIC;
           SAMPLE_OUT : out signed(7 downto 0)
           );
end Tom2;

architecture Behavioral of Tom2 is

type memory is array (0 to 15743) of signed(7 downto 0);
constant tom2_sound: memory := (
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FD",
	x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FE", x"FC", x"FE", x"FC", x"FE", x"FC", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FC", x"FD", x"FC", x"FE", x"FC", x"FE", x"FD", x"FD", x"FD", x"FD", x"FC",
	x"FE", x"FC", x"FF", x"F4", x"B6", x"9E", x"A6", x"A7", x"AE", x"AE", x"BE", x"C1",
	x"CC", x"C8", x"C6", x"D9", x"D7", x"BF", x"E0", x"06", x"FD", x"2C", x"33", x"2E",
	x"20", x"29", x"3B", x"3B", x"35", x"35", x"3D", x"38", x"50", x"6B", x"5E", x"5B",
	x"5F", x"40", x"45", x"4D", x"44", x"2D", x"41", x"38", x"F2", x"17", x"FC", x"EE",
	x"0D", x"C9", x"C1", x"C5", x"AA", x"B4", x"AD", x"9F", x"AE", x"A8", x"AD", x"C4",
	x"B9", x"B8", x"B6", x"B8", x"B3", x"BB", x"CA", x"B5", x"B0", x"BF", x"BF", x"B6",
	x"C6", x"C5", x"CE", x"DD", x"DC", x"B7", x"CA", x"C7", x"B7", x"D3", x"C5", x"CD",
	x"C8", x"EF", x"F6", x"08", x"05", x"0C", x"2D", x"32", x"56", x"6C", x"70", x"63",
	x"68", x"6E", x"6E", x"65", x"61", x"50", x"51", x"57", x"3C", x"41", x"3F", x"40",
	x"43", x"4D", x"3C", x"36", x"31", x"12", x"16", x"E7", x"C8", x"BF", x"C8", x"B5",
	x"AA", x"A4", x"A9", x"C2", x"BE", x"BF", x"BF", x"BE", x"B8", x"9D", x"A5", x"AC",
	x"8F", x"91", x"97", x"B1", x"B4", x"BB", x"BA", x"CD", x"E4", x"E1", x"F0", x"03",
	x"13", x"17", x"37", x"3F", x"45", x"45", x"58", x"62", x"5B", x"6A", x"5B", x"53",
	x"5C", x"65", x"5A", x"52", x"56", x"4F", x"44", x"25", x"2B", x"31", x"41", x"63",
	x"52", x"56", x"56", x"4B", x"4C", x"34", x"40", x"46", x"1E", x"06", x"09", x"0B",
	x"17", x"03", x"EC", x"E1", x"C3", x"BD", x"BE", x"AE", x"A0", x"9C", x"90", x"94",
	x"8B", x"93", x"A6", x"A5", x"96", x"9D", x"9A", x"92", x"99", x"9A", x"99", x"A1",
	x"A0", x"AD", x"CB", x"CD", x"DD", x"F6", x"0F", x"1F", x"35", x"52", x"5F", x"6D",
	x"6F", x"6D", x"70", x"5E", x"65", x"6D", x"62", x"59", x"58", x"62", x"54", x"52",
	x"56", x"5B", x"69", x"6A", x"69", x"61", x"5A", x"47", x"2F", x"25", x"0C", x"08",
	x"FB", x"E4", x"D0", x"BC", x"C1", x"B6", x"AC", x"99", x"96", x"9F", x"8E", x"90",
	x"A3", x"96", x"8C", x"94", x"96", x"99", x"A8", x"AF", x"AA", x"A9", x"AB", x"B8",
	x"C8", x"BE", x"BA", x"BE", x"C6", x"DC", x"E0", x"D0", x"E0", x"EA", x"EC", x"E7",
	x"F9", x"08", x"02", x"17", x"2E", x"40", x"43", x"51", x"57", x"5E", x"66", x"65",
	x"6A", x"6A", x"6D", x"6F", x"73", x"70", x"70", x"71", x"6C", x"6F", x"68", x"6A",
	x"64", x"5A", x"4A", x"46", x"4B", x"37", x"19", x"07", x"F9", x"DB", x"CF", x"B5",
	x"B2", x"A5", x"93", x"8D", x"8C", x"94", x"90", x"90", x"8F", x"8C", x"90", x"92",
	x"8C", x"8D", x"92", x"94", x"8F", x"8D", x"94", x"A0", x"A0", x"99", x"AF", x"C2",
	x"CF", x"E2", x"F1", x"F9", x"F8", x"08", x"23", x"42", x"5A", x"6C", x"73", x"71",
	x"6D", x"62", x"67", x"6F", x"73", x"67", x"63", x"5C", x"56", x"68", x"5D", x"59",
	x"55", x"54", x"59", x"55", x"4B", x"4B", x"4C", x"43", x"30", x"31", x"2E", x"1D",
	x"0F", x"0B", x"0E", x"FD", x"EB", x"DC", x"DA", x"CB", x"BC", x"B4", x"B0", x"A8",
	x"A1", x"A2", x"95", x"93", x"92", x"92", x"90", x"8F", x"97", x"94", x"93", x"91",
	x"8B", x"8F", x"8E", x"8C", x"95", x"96", x"9D", x"A7", x"B6", x"CC", x"E3", x"FC",
	x"0A", x"22", x"39", x"3B", x"38", x"4B", x"55", x"58", x"6C", x"6E", x"70", x"6D",
	x"67", x"71", x"6A", x"68", x"65", x"68", x"6A", x"65", x"6D", x"70", x"6D", x"67",
	x"6A", x"5D", x"4B", x"3F", x"37", x"34", x"1F", x"18", x"08", x"F1", x"E1", x"CD",
	x"B6", x"A6", x"9C", x"93", x"8F", x"8C", x"8F", x"8F", x"8E", x"8C", x"93", x"97",
	x"9A", x"96", x"9D", x"9E", x"95", x"9A", x"9D", x"A2", x"AB", x"B1", x"AB", x"B5",
	x"C3", x"D1", x"DA", x"EB", x"00", x"00", x"09", x"09", x"09", x"11", x"1B", x"21",
	x"27", x"28", x"2D", x"38", x"38", x"46", x"55", x"5D", x"68", x"6E", x"6E", x"72",
	x"72", x"72", x"72", x"71", x"6F", x"74", x"71", x"71", x"6E", x"70", x"60", x"53",
	x"48", x"38", x"28", x"0D", x"F6", x"EB", x"EC", x"E1", x"DA", x"D0", x"C3", x"B5",
	x"A3", x"9B", x"97", x"92", x"92", x"92", x"8E", x"8E", x"8D", x"8C", x"8C", x"8F",
	x"8E", x"8B", x"8D", x"8D", x"92", x"9C", x"AF", x"B9", x"B9", x"BD", x"C4", x"D2",
	x"E2", x"F0", x"F1", x"FE", x"13", x"1A", x"2A", x"41", x"51", x"62", x"69", x"6B",
	x"6E", x"6E", x"6B", x"6A", x"6F", x"6C", x"6A", x"6B", x"6C", x"69", x"69", x"65",
	x"63", x"61", x"61", x"55", x"48", x"3D", x"33", x"2E", x"2C", x"27", x"1E", x"19",
	x"08", x"F8", x"F3", x"EE", x"F0", x"E9", x"DD", x"D1", x"CD", x"C4", x"BA", x"AF",
	x"A8", x"9F", x"9F", x"9D", x"98", x"91", x"91", x"8D", x"8C", x"92", x"92", x"94",
	x"96", x"98", x"96", x"91", x"9D", x"A3", x"AF", x"C4", x"D3", x"E1", x"EF", x"FD",
	x"0B", x"22", x"2B", x"2D", x"30", x"30", x"3F", x"4F", x"59", x"64", x"70", x"71",
	x"71", x"70", x"70", x"6D", x"6B", x"6F", x"72", x"71", x"69", x"63", x"65", x"66",
	x"5E", x"59", x"52", x"4C", x"44", x"38", x"37", x"28", x"14", x"0C", x"FF", x"EE",
	x"E9", x"E2", x"D4", x"C7", x"C2", x"B9", x"B7", x"AD", x"A4", x"9B", x"A0", x"A6",
	x"9E", x"9C", x"9B", x"92", x"93", x"92", x"90", x"98", x"9E", x"A7", x"A4", x"AA",
	x"B6", x"C5", x"C3", x"C3", x"C5", x"CE", x"D0", x"DA", x"E3", x"EB", x"FF", x"00",
	x"00", x"04", x"0D", x"15", x"20", x"2C", x"39", x"49", x"50", x"59", x"5A", x"58",
	x"5D", x"61", x"69", x"70", x"72", x"73", x"73", x"6E", x"6A", x"69", x"69", x"6C",
	x"72", x"66", x"50", x"45", x"36", x"2B", x"21", x"15", x"06", x"FE", x"F8", x"EE",
	x"E0", x"D4", x"C5", x"B5", x"AD", x"A3", x"9E", x"98", x"97", x"90", x"90", x"8F",
	x"8F", x"91", x"97", x"99", x"9F", x"A0", x"A5", x"A8", x"AA", x"B4", x"BA", x"C0",
	x"C3", x"C7", x"CB", x"D9", x"E2", x"EA", x"EB", x"E8", x"E9", x"F4", x"F9", x"03",
	x"0C", x"16", x"21", x"29", x"31", x"32", x"37", x"3E", x"48", x"50", x"5D", x"69",
	x"6C", x"6E", x"6E", x"6A", x"66", x"65", x"5F", x"59", x"5F", x"5F", x"5D", x"5B",
	x"55", x"4A", x"3F", x"38", x"31", x"28", x"24", x"1F", x"1C", x"0E", x"FF", x"F3",
	x"E9", x"E4", x"D7", x"CF", x"C3", x"BD", x"B9", x"AB", x"A0", x"97", x"91", x"94",
	x"90", x"90", x"91", x"8F", x"93", x"92", x"94", x"93", x"97", x"9A", x"9E", x"A3",
	x"A8", x"AE", x"B3", x"BB", x"C2", x"D1", x"E1", x"EF", x"FF", x"07", x"18", x"25",
	x"37", x"42", x"4C", x"54", x"5C", x"64", x"69", x"6A", x"65", x"64", x"60", x"5A",
	x"5B", x"5B", x"5C", x"62", x"5D", x"5B", x"53", x"50", x"4A", x"40", x"3C", x"35",
	x"2F", x"28", x"24", x"1E", x"1A", x"11", x"0C", x"04", x"04", x"FF", x"F7", x"F4",
	x"F2", x"EB", x"E0", x"D8", x"CB", x"C5", x"BD", x"B5", x"AE", x"AC", x"A8", x"A2",
	x"9E", x"A0", x"9E", x"98", x"95", x"94", x"94", x"93", x"97", x"9A", x"A1", x"AC",
	x"B3", x"B9", x"C2", x"CA", x"DA", x"E6", x"EC", x"EF", x"F6", x"FE", x"0B", x"10",
	x"1A", x"22", x"28", x"34", x"3D", x"4A", x"53", x"61", x"67", x"6B", x"6D", x"6A",
	x"6C", x"6B", x"6D", x"6C", x"6E", x"70", x"71", x"70", x"69", x"66", x"61", x"57",
	x"4F", x"41", x"35", x"29", x"19", x"0D", x"04", x"FC", x"F1", x"E7", x"DF", x"D4",
	x"D0", x"C3", x"B6", x"AA", x"A1", x"99", x"97", x"92", x"92", x"92", x"92", x"91",
	x"95", x"97", x"99", x"9F", x"A7", x"AF", x"B4", x"B9", x"BE", x"C4", x"C6", x"C8",
	x"CC", x"D6", x"DF", x"E7", x"EB", x"F1", x"FA", x"01", x"03", x"09", x"10", x"19",
	x"23", x"2A", x"31", x"37", x"3D", x"40", x"45", x"4C", x"51", x"56", x"5D", x"63",
	x"64", x"66", x"68", x"6A", x"67", x"60", x"59", x"5B", x"5A", x"57", x"4F", x"4C",
	x"49", x"44", x"3B", x"31", x"26", x"1E", x"14", x"0C", x"01", x"F5", x"EA", x"DB",
	x"CF", x"C6", x"BD", x"B6", x"AC", x"A1", x"9B", x"95", x"96", x"95", x"91", x"91",
	x"8D", x"8D", x"8B", x"8F", x"93", x"97", x"9F", x"A6", x"AD", x"B2", x"B6", x"BD",
	x"C5", x"CA", x"CF", x"D9", x"E1", x"EE", x"FA", x"06", x"12", x"1C", x"25", x"29",
	x"32", x"3D", x"44", x"4F", x"55", x"5D", x"63", x"6A", x"6F", x"70", x"70", x"73",
	x"71", x"6F", x"6C", x"66", x"5F", x"5E", x"57", x"4F", x"4A", x"44", x"40", x"3A",
	x"30", x"23", x"19", x"15", x"0D", x"00", x"F0", x"E8", x"DE", x"DB", x"D5", x"D0",
	x"CC", x"C6", x"C6", x"C2", x"BF", x"B8", x"B3", x"AE", x"AA", x"A4", x"A0", x"9F",
	x"A0", x"A0", x"A2", x"A5", x"A8", x"AB", x"A8", x"A8", x"A7", x"AC", x"B0", x"B8",
	x"BF", x"C7", x"CE", x"D4", x"DC", x"E4", x"F0", x"FB", x"08", x"15", x"1E", x"2B",
	x"32", x"3B", x"41", x"49", x"4C", x"55", x"5E", x"61", x"67", x"69", x"70", x"73",
	x"73", x"6F", x"6F", x"70", x"6C", x"64", x"59", x"50", x"48", x"42", x"3A", x"34",
	x"33", x"2E", x"28", x"1C", x"15", x"0A", x"01", x"F4", x"E8", x"DE", x"D3", x"CE",
	x"C7", x"C1", x"BA", x"B2", x"AE", x"AB", x"A8", x"A4", x"A0", x"9A", x"97", x"92",
	x"91", x"93", x"92", x"93", x"99", x"9D", x"A5", x"AD", x"B6", x"BE", x"C5", x"CC",
	x"D5", x"DD", x"E5", x"ED", x"F5", x"FE", x"09", x"11", x"1C", x"26", x"27", x"2C",
	x"30", x"32", x"3A", x"41", x"47", x"4C", x"4F", x"50", x"53", x"55", x"56", x"5B",
	x"5B", x"5B", x"59", x"58", x"55", x"53", x"53", x"4F", x"4D", x"46", x"41", x"3B",
	x"34", x"2C", x"24", x"1C", x"16", x"0F", x"0A", x"05", x"FE", x"F5", x"E9", x"DE",
	x"D2", x"CA", x"C2", x"BE", x"B4", x"B1", x"AB", x"A8", x"A4", x"9D", x"9B", x"98",
	x"97", x"96", x"9A", x"9C", x"A0", x"A5", x"AA", x"AE", x"B1", x"BC", x"C4", x"CD",
	x"D5", x"DA", x"E3", x"EA", x"F3", x"F8", x"FF", x"04", x"0C", x"14", x"1F", x"25",
	x"2D", x"32", x"37", x"3C", x"3D", x"43", x"45", x"49", x"4C", x"50", x"53", x"54",
	x"57", x"56", x"58", x"57", x"56", x"52", x"4E", x"49", x"47", x"44", x"3F", x"39",
	x"30", x"2B", x"24", x"1D", x"13", x"0C", x"03", x"FC", x"F5", x"EF", x"E9", x"E4",
	x"DD", x"D6", x"D1", x"CA", x"C6", x"C0", x"BB", x"B4", x"B2", x"AF", x"AF", x"AD",
	x"AF", x"AF", x"B0", x"B0", x"B1", x"B2", x"B6", x"B8", x"BE", x"C2", x"C6", x"C9",
	x"CF", x"D4", x"D9", x"DF", x"E4", x"E8", x"ED", x"F2", x"F6", x"FD", x"03", x"09",
	x"11", x"18", x"1F", x"29", x"30", x"36", x"3D", x"41", x"45", x"49", x"4B", x"4F",
	x"50", x"55", x"57", x"57", x"56", x"55", x"50", x"4E", x"4A", x"48", x"45", x"3E",
	x"3A", x"30", x"29", x"1F", x"18", x"14", x"0E", x"0A", x"01", x"FA", x"F2", x"EC",
	x"E6", x"E1", x"DB", x"D5", x"D2", x"CD", x"CA", x"C8", x"C7", x"C3", x"C1", x"BD",
	x"BA", x"BB", x"BA", x"BC", x"BD", x"C0", x"BF", x"BD", x"BB", x"BA", x"BD", x"C0",
	x"C1", x"C5", x"C8", x"CF", x"D1", x"D6", x"DC", x"E1", x"E9", x"EF", x"F7", x"FD",
	x"04", x"0A", x"12", x"18", x"20", x"27", x"2D", x"33", x"3A", x"3F", x"47", x"4C",
	x"4E", x"4F", x"4C", x"4A", x"47", x"47", x"45", x"45", x"44", x"42", x"41", x"40",
	x"3E", x"3B", x"38", x"35", x"2D", x"26", x"20", x"19", x"12", x"0C", x"05", x"00",
	x"FB", x"F5", x"F1", x"ED", x"E8", x"E5", x"E1", x"DA", x"D8", x"D1", x"CC", x"C7",
	x"C2", x"BE", x"BC", x"B7", x"B4", x"B2", x"AF", x"AF", x"B0", x"B3", x"B3", x"B8",
	x"BC", x"BF", x"C4", x"C7", x"CA", x"CF", x"D3", x"DC", x"E3", x"EB", x"F2", x"F9",
	x"00", x"06", x"0D", x"11", x"17", x"19", x"1B", x"22", x"24", x"28", x"2A", x"2E",
	x"33", x"35", x"3B", x"3E", x"43", x"44", x"46", x"46", x"45", x"46", x"44", x"46",
	x"44", x"44", x"43", x"3E", x"39", x"35", x"30", x"2D", x"27", x"23", x"1D", x"18",
	x"13", x"0D", x"07", x"00", x"FB", x"F6", x"EF", x"E8", x"E1", x"DB", x"D3", x"CE",
	x"C7", x"C0", x"BB", x"B7", x"B2", x"B0", x"AD", x"AD", x"AC", x"AE", x"AF", x"B2",
	x"B5", x"B8", x"BE", x"C2", x"C9", x"CC", x"D2", x"D4", x"D9", x"DD", x"E3", x"E7",
	x"EC", x"F1", x"F7", x"FB", x"02", x"07", x"0D", x"12", x"17", x"1E", x"21", x"26",
	x"2C", x"32", x"37", x"3C", x"3E", x"42", x"42", x"45", x"45", x"47", x"48", x"47",
	x"49", x"47", x"49", x"48", x"45", x"43", x"3E", x"39", x"34", x"2F", x"29", x"25",
	x"20", x"1C", x"14", x"0F", x"05", x"FE", x"F7", x"EE", x"E7", x"E0", x"D9", x"D4",
	x"CE", x"CB", x"C6", x"C3", x"BF", x"B9", x"B7", x"B3", x"B3", x"B1", x"B3", x"B3",
	x"B6", x"B7", x"BB", x"BF", x"C2", x"C7", x"C9", x"CD", x"D0", x"D3", x"D4", x"D8",
	x"D9", x"DF", x"E4", x"E8", x"F0", x"F6", x"FD", x"01", x"07", x"0C", x"10", x"17",
	x"1B", x"23", x"2A", x"30", x"39", x"3E", x"46", x"4A", x"50", x"52", x"52", x"54",
	x"51", x"51", x"4E", x"4C", x"48", x"45", x"42", x"41", x"3E", x"3C", x"36", x"2E",
	x"29", x"21", x"1A", x"10", x"09", x"01", x"FC", x"F6", x"F0", x"EC", x"E5", x"E0",
	x"DB", x"D6", x"D4", x"CF", x"CD", x"CB", x"C8", x"C5", x"C2", x"BE", x"BA", x"B9",
	x"B6", x"B6", x"B5", x"B7", x"B6", x"B8", x"B8", x"BB", x"BB", x"BF", x"C1", x"C5",
	x"C9", x"CF", x"D5", x"DC", x"E4", x"EB", x"F2", x"FB", x"03", x"0A", x"12", x"18",
	x"1F", x"25", x"2A", x"2F", x"34", x"39", x"40", x"45", x"48", x"4C", x"4C", x"4E",
	x"4D", x"4E", x"4D", x"4C", x"4B", x"45", x"43", x"3D", x"37", x"34", x"30", x"2C",
	x"29", x"24", x"1F", x"19", x"15", x"0E", x"0A", x"05", x"01", x"FA", x"F6", x"F1",
	x"EE", x"EA", x"E5", x"E0", x"DA", x"D3", x"CF", x"CA", x"C8", x"C5", x"C4", x"C1",
	x"BF", x"BC", x"BB", x"B7", x"B8", x"B7", x"B5", x"B7", x"B8", x"BC", x"BF", x"C4",
	x"C8", x"CE", x"D2", x"D9", x"DD", x"E0", x"E6", x"E9", x"F0", x"F5", x"FC", x"03",
	x"08", x"0F", x"16", x"1C", x"22", x"29", x"2D", x"33", x"37", x"3C", x"40", x"43",
	x"45", x"45", x"46", x"47", x"46", x"47", x"47", x"48", x"47", x"47", x"45", x"43",
	x"3E", x"38", x"32", x"2C", x"26", x"20", x"19", x"16", x"12", x"0F", x"0A", x"05",
	x"FE", x"F8", x"F0", x"EA", x"E2", x"DC", x"D4", x"CF", x"C9", x"C5", x"C1", x"BB",
	x"B8", x"B4", x"B3", x"B2", x"B0", x"B1", x"B2", x"B4", x"B5", x"B8", x"BA", x"C0",
	x"C3", x"C9", x"CE", x"D5", x"DB", x"E0", x"E7", x"EB", x"F2", x"F6", x"FB", x"00",
	x"04", x"0B", x"0E", x"14", x"17", x"1C", x"20", x"23", x"25", x"28", x"29", x"2C",
	x"2E", x"32", x"35", x"38", x"3B", x"3D", x"3D", x"3E", x"3E", x"3E", x"3C", x"3D",
	x"3B", x"3B", x"3A", x"3A", x"38", x"36", x"31", x"2D", x"29", x"24", x"20", x"1A",
	x"14", x"0D", x"05", x"FD", x"F6", x"ED", x"E7", x"DF", x"DA", x"D3", x"CF", x"CA",
	x"C7", x"C2", x"C0", x"BD", x"BC", x"B9", x"B8", x"B5", x"B5", x"B3", x"B5", x"B5",
	x"B9", x"BB", x"C0", x"C4", x"C6", x"CC", x"CF", x"D4", x"D7", x"DB", x"DF", x"E4",
	x"EA", x"F0", x"F8", x"FF", x"06", x"0C", x"10", x"16", x"1A", x"1F", x"24", x"27",
	x"2D", x"32", x"38", x"3D", x"40", x"46", x"49", x"4F", x"51", x"53", x"52", x"52",
	x"4E", x"4C", x"47", x"43", x"3E", x"3A", x"33", x"2F", x"28", x"23", x"1C", x"18",
	x"11", x"0C", x"03", x"FD", x"F5", x"EF", x"E8", x"E5", x"E0", x"DC", x"DA", x"D6",
	x"D2", x"D0", x"CB", x"C9", x"C6", x"C4", x"C1", x"C2", x"C0", x"C1", x"C1", x"C3",
	x"C3", x"C6", x"C5", x"C7", x"C6", x"C8", x"C8", x"CA", x"CA", x"CE", x"D2", x"D6",
	x"DA", x"DD", x"E3", x"E9", x"EF", x"F3", x"FA", x"FF", x"06", x"0B", x"13", x"19",
	x"1F", x"27", x"2C", x"33", x"38", x"3F", x"42", x"44", x"48", x"47", x"49", x"49",
	x"4A", x"49", x"4B", x"4A", x"4A", x"47", x"46", x"41", x"3F", x"3B", x"36", x"30",
	x"2A", x"22", x"1C", x"13", x"0D", x"05", x"00", x"FA", x"F3", x"F0", x"EA", x"E6",
	x"E1", x"D9", x"D4", x"CD", x"C9", x"C4", x"C0", x"BD", x"B9", x"B6", x"B4", x"B2",
	x"B2", x"B1", x"B2", x"B2", x"B5", x"B7", x"BB", x"BC", x"C0", x"C2", x"C6", x"CB",
	x"CF", x"D7", x"DD", x"E6", x"ED", x"F3", x"FB", x"00", x"08", x"0D", x"13", x"17",
	x"1E", x"22", x"29", x"2E", x"35", x"3A", x"41", x"45", x"49", x"4A", x"4B", x"48",
	x"48", x"46", x"44", x"41", x"3E", x"3E", x"3B", x"39", x"35", x"34", x"30", x"2C",
	x"29", x"24", x"21", x"1D", x"19", x"14", x"0F", x"0C", x"06", x"02", x"FB", x"F8",
	x"F3", x"EE", x"E9", x"E2", x"DE", x"D9", x"D2", x"CE", x"C8", x"C4", x"BF", x"B9",
	x"B7", x"B4", x"B1", x"B0", x"AF", x"B0", x"B0", x"B1", x"B4", x"B8", x"BC", x"C0",
	x"C6", x"CC", x"CF", x"D6", x"DB", x"E1", x"E7", x"EE", x"F3", x"FA", x"FF", x"06",
	x"0D", x"13", x"1A", x"21", x"28", x"2E", x"33", x"37", x"3B", x"3F", x"42", x"47",
	x"4A", x"4A", x"4C", x"4B", x"4D", x"4B", x"4A", x"49", x"46", x"45", x"41", x"3C",
	x"38", x"33", x"2E", x"28", x"24", x"1E", x"1A", x"16", x"0F", x"0B", x"05", x"00",
	x"F8", x"F2", x"EA", x"E4", x"DB", x"D5", x"CE", x"C7", x"C3", x"BD", x"BB", x"B9",
	x"B5", x"B4", x"B2", x"B2", x"B2", x"B1", x"B4", x"B7", x"BB", x"BF", x"C5", x"CA",
	x"CD", x"D2", x"D6", x"DA", x"DD", x"E3", x"E7", x"ED", x"F1", x"F7", x"FB", x"00",
	x"04", x"09", x"0C", x"10", x"14", x"18", x"1D", x"22", x"26", x"2A", x"2C", x"30",
	x"33", x"34", x"38", x"3A", x"3D", x"3F", x"40", x"43", x"45", x"44", x"46", x"44",
	x"43", x"41", x"3D", x"3B", x"35", x"31", x"2B", x"26", x"20", x"1A", x"13", x"0D",
	x"06", x"FF", x"F7", x"F1", x"EA", x"E5", x"E0", x"DB", x"D7", x"D4", x"D0", x"CE",
	x"CA", x"C6", x"C5", x"C1", x"BF", x"BD", x"BA", x"B8", x"B6", x"B7", x"B7", x"BB",
	x"BE", x"C1", x"C6", x"C9", x"CC", x"D1", x"D3", x"D8", x"DB", x"E0", x"E5", x"EA",
	x"F1", x"F6", x"FE", x"04", x"0B", x"10", x"17", x"1B", x"1D", x"22", x"25", x"28",
	x"2C", x"30", x"36", x"3A", x"3E", x"43", x"44", x"47", x"46", x"47", x"46", x"45",
	x"44", x"40", x"3F", x"3D", x"38", x"35", x"2F", x"2A", x"23", x"1F", x"1A", x"14",
	x"10", x"0A", x"03", x"FE", x"F6", x"F1", x"EA", x"E6", x"E1", x"DC", x"DA", x"D7",
	x"D4", x"D3", x"D1", x"D1", x"D0", x"CF", x"CD", x"CA", x"C9", x"C7", x"C7", x"C5",
	x"C6", x"C7", x"C7", x"C9", x"C9", x"CC", x"CD", x"CF", x"D2", x"D4", x"D8", x"DB",
	x"DE", x"E3", x"E8", x"EC", x"F2", x"F7", x"FC", x"01", x"07", x"0D", x"11", x"17",
	x"1B", x"21", x"25", x"29", x"2D", x"32", x"35", x"3A", x"3C", x"3D", x"40", x"3F",
	x"41", x"41", x"40", x"41", x"3F", x"3F", x"3D", x"3A", x"35", x"32", x"2C", x"28",
	x"21", x"1D", x"18", x"13", x"0D", x"0A", x"05", x"02", x"FD", x"F9", x"F4", x"F0",
	x"EB", x"E6", x"DF", x"DB", x"D5", x"D1", x"CC", x"C9", x"C6", x"C4", x"C1", x"BF",
	x"C0", x"BE", x"BF", x"BF", x"C0", x"C0", x"C2", x"C3", x"C4", x"C7", x"C9", x"CE",
	x"D0", x"D5", x"D9", x"DF", x"E4", x"E9", x"F1", x"F7", x"FC", x"04", x"08", x"0F",
	x"13", x"19", x"1E", x"23", x"29", x"2D", x"33", x"37", x"3A", x"3B", x"3D", x"3C",
	x"3B", x"3A", x"37", x"37", x"34", x"34", x"33", x"31", x"31", x"2E", x"2D", x"2B",
	x"29", x"26", x"23", x"1F", x"1C", x"18", x"15", x"11", x"0D", x"0A", x"06", x"04",
	x"FF", x"FC", x"F6", x"F2", x"EC", x"E8", x"E2", x"DE", x"D9", x"D4", x"D0", x"CC",
	x"C9", x"C4", x"C2", x"BF", x"BD", x"BC", x"BE", x"BE", x"C0", x"C1", x"C4", x"C6",
	x"C9", x"CC", x"CF", x"D4", x"D7", x"DC", x"E0", x"E3", x"E9", x"ED", x"F1", x"F7",
	x"FB", x"01", x"06", x"09", x"0F", x"12", x"18", x"1C", x"22", x"26", x"2C", x"2F",
	x"35", x"38", x"3A", x"3D", x"3E", x"3D", x"3F", x"3F", x"40", x"40", x"3E", x"3E",
	x"3C", x"3A", x"37", x"34", x"2F", x"2C", x"28", x"23", x"1F", x"19", x"15", x"0E",
	x"0A", x"04", x"FE", x"F9", x"F4", x"EE", x"E9", x"E3", x"DC", x"D7", x"D2", x"CC",
	x"C9", x"C6", x"C5", x"C3", x"C1", x"C0", x"BF", x"C0", x"C0", x"C2", x"C2", x"C5",
	x"C6", x"C9", x"CB", x"CF", x"D1", x"D6", x"DA", x"DD", x"E3", x"E7", x"EC", x"EF",
	x"F4", x"F7", x"FC", x"FF", x"04", x"08", x"0B", x"0E", x"12", x"16", x"19", x"1D",
	x"20", x"23", x"26", x"2A", x"2D", x"30", x"32", x"36", x"37", x"3A", x"3A", x"3C",
	x"3B", x"3C", x"3C", x"3A", x"3A", x"37", x"35", x"31", x"2D", x"29", x"23", x"1F",
	x"19", x"15", x"0F", x"0C", x"06", x"02", x"FD", x"F9", x"F3", x"EE", x"E9", x"E4",
	x"DF", x"D9", x"D5", x"CF", x"CD", x"CA", x"C7", x"C6", x"C3", x"C3", x"C2", x"C2",
	x"C2", x"C3", x"C4", x"C5", x"C8", x"CB", x"CB", x"CE", x"D0", x"D4", x"D7", x"D9",
	x"DF", x"E2", x"E8", x"EC", x"F2", x"F6", x"FC", x"FF", x"04", x"08", x"0D", x"10",
	x"15", x"19", x"1E", x"22", x"27", x"2B", x"30", x"33", x"37", x"38", x"3A", x"3D",
	x"3D", x"3F", x"3E", x"3E", x"3D", x"3B", x"3A", x"37", x"35", x"31", x"2D", x"2A",
	x"25", x"20", x"19", x"15", x"0F", x"0A", x"04", x"00", x"FB", x"F5", x"F1", x"EC",
	x"EA", x"E6", x"E2", x"E0", x"DD", x"DB", x"DA", x"D7", x"D6", x"D5", x"D2", x"D1",
	x"CF", x"CC", x"CC", x"CA", x"CB", x"CA", x"CB", x"CB", x"CD", x"CF", x"D0", x"D1",
	x"D4", x"D6", x"D9", x"DB", x"DF", x"E1", x"E6", x"E9", x"EF", x"F4", x"F8", x"FF",
	x"03", x"08", x"0F", x"12", x"17", x"1B", x"1E", x"23", x"25", x"2A", x"2D", x"32",
	x"35", x"38", x"3A", x"3B", x"3C", x"3B", x"3B", x"38", x"37", x"35", x"33", x"30",
	x"2E", x"2A", x"28", x"24", x"22", x"1D", x"1A", x"15", x"13", x"0E", x"0B", x"07",
	x"04", x"FF", x"FC", x"F6", x"F3", x"EE", x"E8", x"E5", x"E0", x"DD", x"D9", x"D7",
	x"D4", x"D0", x"CE", x"CA", x"C8", x"C5", x"C5", x"C4", x"C3", x"C5", x"C4", x"C6",
	x"C7", x"CB", x"CE", x"D0", x"D4", x"D7", x"DA", x"DE", x"E1", x"E7", x"EB", x"F1",
	x"F5", x"FB", x"01", x"05", x"0B", x"0F", x"14", x"17", x"1C", x"20", x"22", x"26",
	x"28", x"2C", x"2E", x"2F", x"30", x"31", x"32", x"32", x"34", x"33", x"35", x"33",
	x"32", x"31", x"2E", x"2D", x"2A", x"28", x"27", x"25", x"23", x"1F", x"1D", x"19",
	x"14", x"11", x"0D", x"07", x"05", x"FF", x"FC", x"F7", x"F4", x"EF", x"E9", x"E6",
	x"E0", x"DD", x"D8", x"D4", x"D0", x"CE", x"CB", x"CA", x"C8", x"C6", x"C6", x"C5",
	x"C6", x"C6", x"C8", x"CA", x"CA", x"CD", x"CE", x"D2", x"D4", x"D8", x"DC", x"DE",
	x"E3", x"E6", x"EC", x"F0", x"F4", x"FA", x"FE", x"03", x"07", x"0C", x"0F", x"14",
	x"17", x"1C", x"20", x"23", x"28", x"2A", x"2E", x"2F", x"32", x"33", x"33", x"35",
	x"35", x"36", x"36", x"35", x"36", x"34", x"34", x"32", x"31", x"2F", x"2B", x"29",
	x"25", x"22", x"1C", x"19", x"13", x"10", x"0A", x"06", x"FF", x"FB", x"F5", x"F1",
	x"EB", x"E7", x"E3", x"DF", x"DC", x"D7", x"D5", x"D1", x"D0", x"CC", x"CA", x"C7",
	x"C7", x"C6", x"C5", x"C6", x"C6", x"C6", x"C9", x"CA", x"CE", x"CF", x"D4", x"D6",
	x"DA", x"DE", x"E0", x"E5", x"E7", x"EC", x"EF", x"F4", x"F8", x"FB", x"00", x"04",
	x"08", x"0B", x"10", x"12", x"17", x"19", x"1C", x"20", x"23", x"27", x"2A", x"2D",
	x"31", x"33", x"37", x"38", x"39", x"3A", x"39", x"39", x"38", x"37", x"34", x"33",
	x"30", x"2E", x"2B", x"27", x"22", x"1F", x"19", x"16", x"10", x"0C", x"06", x"02",
	x"FC", x"F8", x"F3", x"ED", x"EA", x"E4", x"E0", x"DC", x"D7", x"D5", x"D1", x"D0",
	x"CE", x"CD", x"CC", x"CA", x"CA", x"C9", x"CA", x"C9", x"CB", x"CC", x"CE", x"CF",
	x"D2", x"D3", x"D7", x"D9", x"DB", x"DE", x"E0", x"E4", x"E5", x"E9", x"EC", x"EE",
	x"F3", x"F6", x"FC", x"FF", x"05", x"09", x"10", x"14", x"1A", x"1D", x"23", x"27",
	x"2B", x"2E", x"32", x"34", x"37", x"38", x"3A", x"3A", x"3B", x"3B", x"3A", x"38",
	x"35", x"34", x"30", x"2F", x"2A", x"28", x"23", x"1F", x"1C", x"16", x"13", x"0F",
	x"09", x"06", x"01", x"FE", x"F9", x"F6", x"F2", x"ED", x"EB", x"E6", x"E4", x"DF",
	x"DD", x"DA", x"D6", x"D4", x"D1", x"D0", x"CE", x"CD", x"CB", x"CC", x"CA", x"CB",
	x"CB", x"CA", x"CC", x"CD", x"CD", x"D1", x"D2", x"D6", x"D9", x"DE", x"E1", x"E5",
	x"E8", x"EC", x"F1", x"F4", x"FA", x"FE", x"01", x"07", x"0B", x"0F", x"14", x"18",
	x"1B", x"21", x"24", x"28", x"2A", x"2E", x"2F", x"32", x"32", x"33", x"33", x"33",
	x"33", x"31", x"31", x"30", x"2E", x"2E", x"2B", x"2B", x"28", x"26", x"22", x"20",
	x"1C", x"18", x"13", x"10", x"0C", x"09", x"04", x"01", x"FD", x"F8", x"F5", x"EF",
	x"EC", x"E9", x"E4", x"E2", x"DE", x"DC", x"D9", x"D7", x"D4", x"D2", x"D1", x"CE",
	x"CE", x"CC", x"CA", x"CB", x"C9", x"CA", x"C9", x"CC", x"CD", x"D0", x"D2", x"D7",
	x"DB", x"DF", x"E2", x"E6", x"EB", x"EE", x"F4", x"F8", x"FB", x"01", x"04", x"0A",
	x"0E", x"11", x"15", x"18", x"1C", x"1E", x"22", x"23", x"26", x"28", x"2B", x"2C",
	x"2F", x"30", x"30", x"32", x"31", x"32", x"30", x"30", x"2E", x"2D", x"2B", x"28",
	x"26", x"22", x"20", x"1C", x"1A", x"15", x"13", x"0F", x"0D", x"0A", x"05", x"03",
	x"FE", x"FC", x"F8", x"F3", x"F0", x"EB", x"E8", x"E3", x"E1", x"DC", x"DA", x"D6",
	x"D5", x"D2", x"D1", x"CE", x"CE", x"CD", x"CB", x"CC", x"CB", x"CC", x"CD", x"CF",
	x"D0", x"D3", x"D5", x"D9", x"DD", x"DF", x"E4", x"E6", x"EB", x"EE", x"F3", x"F6",
	x"FB", x"FE", x"04", x"07", x"0C", x"10", x"13", x"17", x"1A", x"1C", x"1F", x"20",
	x"23", x"23", x"26", x"26", x"29", x"2A", x"2B", x"2D", x"2D", x"2E", x"2D", x"2F",
	x"2D", x"2E", x"2D", x"2B", x"2B", x"28", x"26", x"23", x"20", x"1D", x"18", x"15",
	x"10", x"0C", x"08", x"02", x"FF", x"F9", x"F6", x"F2", x"EC", x"E9", x"E4", x"E1",
	x"DC", x"D9", x"D5", x"D4", x"D1", x"D1", x"D0", x"CE", x"CF", x"CF", x"CE", x"D0",
	x"D0", x"D2", x"D3", x"D6", x"D6", x"D9", x"DB", x"DC", x"E0", x"E1", x"E4", x"E7",
	x"E9", x"ED", x"EF", x"F3", x"F5", x"FA", x"FC", x"01", x"04", x"08", x"0C", x"0E",
	x"13", x"16", x"1B", x"1E", x"22", x"26", x"28", x"2C", x"2D", x"30", x"30", x"32",
	x"31", x"32", x"31", x"31", x"2F", x"2F", x"2D", x"2C", x"2A", x"27", x"26", x"21",
	x"1F", x"1B", x"17", x"11", x"0E", x"08", x"05", x"00", x"FD", x"F9", x"F6", x"F1",
	x"EF", x"EA", x"E8", x"E4", x"E0", x"DE", x"DA", x"D8", x"D6", x"D3", x"D3", x"D1",
	x"D1", x"D1", x"D0", x"D1", x"D0", x"D2", x"D2", x"D5", x"D5", x"D7", x"DA", x"DB",
	x"DE", x"E0", x"E1", x"E5", x"E7", x"EB", x"ED", x"F2", x"F5", x"F9", x"FD", x"01",
	x"04", x"08", x"0C", x"10", x"14", x"18", x"1A", x"1F", x"23", x"25", x"2A", x"2C",
	x"2F", x"30", x"32", x"31", x"32", x"31", x"31", x"2F", x"2F", x"2D", x"2A", x"29",
	x"26", x"25", x"21", x"1F", x"1B", x"18", x"14", x"10", x"0D", x"09", x"06", x"02",
	x"00", x"FB", x"F9", x"F4", x"F1", x"EC", x"EA", x"E6", x"E3", x"E0", x"DD", x"DB",
	x"D8", x"D7", x"D4", x"D3", x"D1", x"D1", x"D0", x"CF", x"D0", x"CF", x"D2", x"D2",
	x"D4", x"D6", x"D9", x"DA", x"DD", x"DF", x"E3", x"E5", x"E8", x"EA", x"EE", x"F2",
	x"F4", x"F9", x"FB", x"00", x"03", x"08", x"0C", x"11", x"15", x"19", x"1C", x"1E",
	x"22", x"24", x"27", x"29", x"2A", x"2C", x"2C", x"2E", x"2E", x"2F", x"2E", x"2F",
	x"2D", x"2D", x"2C", x"29", x"27", x"24", x"21", x"1D", x"1B", x"16", x"14", x"0F",
	x"0D", x"0A", x"05", x"03", x"FF", x"FC", x"F9", x"F5", x"F3", x"F0", x"ED", x"EA",
	x"E7", x"E5", x"E2", x"E1", x"DF", x"DD", x"DA", x"D8", x"D5", x"D4", x"D1", x"D0",
	x"CE", x"CE", x"CD", x"CE", x"CE", x"D1", x"D2", x"D6", x"D9", x"DC", x"E0", x"E3",
	x"E7", x"EB", x"F0", x"F4", x"F7", x"FD", x"00", x"05", x"08", x"0C", x"0E", x"12",
	x"14", x"17", x"19", x"1C", x"1D", x"21", x"23", x"24", x"26", x"27", x"28", x"28",
	x"29", x"29", x"2A", x"29", x"2A", x"28", x"29", x"27", x"25", x"25", x"22", x"21",
	x"1F", x"1B", x"19", x"15", x"13", x"0F", x"0D", x"09", x"04", x"01", x"FC", x"F9",
	x"F6", x"F1", x"EE", x"EA", x"E7", x"E4", x"E0", x"DE", x"DB", x"D8", x"D7", x"D5",
	x"D3", x"D3", x"D3", x"D2", x"D1", x"D3", x"D2", x"D4", x"D4", x"D6", x"D8", x"DA",
	x"DC", x"DE", x"E1", x"E4", x"E8", x"EB", x"EE", x"F2", x"F5", x"FA", x"FD", x"00",
	x"04", x"06", x"0A", x"0D", x"0E", x"12", x"15", x"16", x"1A", x"1C", x"1F", x"20",
	x"24", x"26", x"27", x"28", x"29", x"29", x"2B", x"2A", x"2B", x"2A", x"2A", x"29",
	x"28", x"26", x"25", x"22", x"21", x"1D", x"1B", x"17", x"15", x"10", x"0E", x"09",
	x"07", x"02", x"FF", x"FA", x"F7", x"F2", x"EF", x"EB", x"E7", x"E4", x"E1", x"DE",
	x"DC", x"DA", x"D8", x"D5", x"D5", x"D4", x"D5", x"D4", x"D6", x"D6", x"D6", x"D7",
	x"D7", x"D9", x"DA", x"DA", x"DD", x"DF", x"E0", x"E3", x"E5", x"E8", x"EA", x"EE",
	x"F0", x"F3", x"F6", x"F9", x"FD", x"FF", x"04", x"07", x"0C", x"10", x"13", x"17",
	x"1B", x"1D", x"20", x"22", x"25", x"25", x"28", x"29", x"29", x"2A", x"2B", x"2A",
	x"2B", x"2A", x"2A", x"29", x"28", x"27", x"24", x"23", x"20", x"1E", x"1B", x"18",
	x"16", x"12", x"0F", x"0C", x"08", x"05", x"01", x"FC", x"F9", x"F5", x"F0", x"ED",
	x"E9", x"E4", x"E2", x"DF", x"DE", x"DB", x"DA", x"D8", x"D7", x"D6", x"D4", x"D5",
	x"D4", x"D5", x"D5", x"D5", x"D7", x"D8", x"DA", x"DB", x"DD", x"DE", x"E1", x"E2",
	x"E5", x"E8", x"E9", x"ED", x"F0", x"F1", x"F5", x"F7", x"FB", x"FE", x"00", x"04",
	x"07", x"0B", x"0F", x"11", x"16", x"19", x"1D", x"20", x"24", x"26", x"2A", x"2B",
	x"2E", x"2E", x"2F", x"2F", x"2F", x"2E", x"2D", x"2B", x"2A", x"27", x"25", x"21",
	x"1F", x"1C", x"18", x"16", x"12", x"0F", x"0C", x"08", x"06", x"03", x"FF", x"FD",
	x"FA", x"F6", x"F4", x"F2", x"EE", x"EC", x"E8", x"E6", x"E4", x"E0", x"DF", x"DC",
	x"DB", x"D9", x"D7", x"D7", x"D5", x"D5", x"D4", x"D4", x"D5", x"D4", x"D6", x"D6",
	x"D9", x"DA", x"DC", x"DE", x"E1", x"E2", x"E6", x"E9", x"ED", x"F1", x"F4", x"F9",
	x"FC", x"01", x"05", x"08", x"0C", x"0F", x"12", x"15", x"18", x"1B", x"1D", x"1F",
	x"22", x"23", x"26", x"27", x"29", x"2A", x"2B", x"2B", x"29", x"2A", x"28", x"28",
	x"26", x"26", x"23", x"22", x"1F", x"1E", x"1A", x"18", x"14", x"12", x"0E", x"0A",
	x"08", x"04", x"02", x"FE", x"FC", x"F9", x"F7", x"F3", x"F2", x"EF", x"EB", x"EA",
	x"E6", x"E4", x"E0", x"DE", x"DC", x"D8", x"D8", x"D5", x"D5", x"D4", x"D4", x"D3",
	x"D4", x"D4", x"D5", x"D7", x"D7", x"DA", x"DC", x"DD", x"E1", x"E4", x"E7", x"EB",
	x"EE", x"F2", x"F6", x"F9", x"FD", x"FF", x"04", x"06", x"0A", x"0D", x"0F", x"13",
	x"15", x"18", x"1A", x"1B", x"1D", x"1F", x"20", x"22", x"22", x"24", x"24", x"26",
	x"27", x"26", x"27", x"26", x"27", x"26", x"24", x"24", x"22", x"1F", x"1E", x"1B",
	x"19", x"16", x"14", x"10", x"0D", x"09", x"06", x"02", x"FF", x"FA", x"F8", x"F4",
	x"F1", x"EE", x"EB", x"E7", x"E6", x"E4", x"E1", x"E0", x"DD", x"DC", x"DA", x"D9",
	x"D7", x"D7", x"D6", x"D5", x"D6", x"D5", x"D6", x"D8", x"D8", x"DB", x"DC", x"DF",
	x"E1", x"E4", x"E7", x"E9", x"ED", x"EF", x"F4", x"F6", x"FA", x"FD", x"01", x"03",
	x"07", x"09", x"0D", x"10", x"12", x"15", x"17", x"1A", x"1B", x"1E", x"1E", x"21",
	x"22", x"22", x"24", x"23", x"25", x"24", x"25", x"24", x"25", x"24", x"22", x"22",
	x"21", x"1E", x"1E", x"1B", x"1A", x"19", x"15", x"14", x"11", x"0E", x"0B", x"07",
	x"04", x"00", x"FD", x"F8", x"F5", x"F1", x"EE", x"EA", x"E8", x"E4", x"E2", x"DF",
	x"DE", x"DC", x"DA", x"D9", x"D8", x"D8", x"D8", x"D8", x"D8", x"D9", x"D9", x"DB",
	x"DB", x"DE", x"DF", x"E2", x"E3", x"E6", x"E8", x"E9", x"EB", x"ED", x"EF", x"F2",
	x"F5", x"F8", x"FB", x"FE", x"00", x"03", x"05", x"09", x"0B", x"0F", x"11", x"15",
	x"17", x"1B", x"1D", x"1F", x"22", x"23", x"26", x"27", x"27", x"28", x"27", x"28",
	x"27", x"27", x"25", x"25", x"23", x"23", x"20", x"1F", x"1D", x"19", x"17", x"13",
	x"10", x"0C", x"09", x"05", x"02", x"FE", x"FB", x"F7", x"F5", x"F1", x"EF", x"EB",
	x"EA", x"E7", x"E4", x"E3", x"E0", x"DF", x"DE", x"DD", x"DC", x"DB", x"DB", x"DA",
	x"DB", x"DA", x"DC", x"DC", x"DD", x"DE", x"DE", x"E0", x"E1", x"E3", x"E5", x"E5",
	x"E8", x"EA", x"ED", x"EE", x"F2", x"F3", x"F7", x"F9", x"FD", x"FF", x"03", x"06",
	x"08", x"0D", x"0F", x"13", x"15", x"19", x"1C", x"1E", x"21", x"22", x"25", x"25",
	x"27", x"27", x"28", x"27", x"28", x"26", x"26", x"23", x"23", x"21", x"1E", x"1D",
	x"1A", x"19", x"15", x"14", x"10", x"0F", x"0B", x"09", x"05", x"03", x"FF", x"FD",
	x"F9", x"F7", x"F3", x"F2", x"EE", x"ED", x"EA", x"E8", x"E6", x"E4", x"E1", x"E0",
	x"DD", x"DD", x"DC", x"DA", x"DA", x"D8", x"D9", x"D8", x"D9", x"D8", x"DA", x"DB",
	x"DC", x"DE", x"E0", x"E2", x"E5", x"E8", x"EA", x"EE", x"F0", x"F5", x"F8", x"FA",
	x"FE", x"00", x"04", x"07", x"0B", x"0D", x"0F", x"13", x"15", x"18", x"19", x"1C",
	x"1E", x"1F", x"21", x"23", x"23", x"25", x"25", x"27", x"26", x"27", x"25", x"25",
	x"24", x"21", x"20", x"1D", x"1B", x"18", x"17", x"13", x"12", x"0F", x"0C", x"0A",
	x"07", x"04", x"02", x"FE", x"FD", x"F9", x"F7", x"F4", x"F1", x"EF", x"EC", x"EB",
	x"E9", x"E6", x"E5", x"E2", x"E1", x"DE", x"DE", x"DB", x"DB", x"DA", x"DA", x"DA",
	x"D9", x"DB", x"DA", x"DC", x"DD", x"DF", x"DF", x"E2", x"E4", x"E6", x"E9", x"EB",
	x"ED", x"F1", x"F4", x"F8", x"FB", x"FE", x"01", x"05", x"07", x"0B", x"0D", x"11",
	x"13", x"16", x"17", x"1A", x"1B", x"1D", x"1F", x"20", x"21", x"22", x"21", x"22",
	x"23", x"23", x"23", x"22", x"21", x"21", x"1F", x"1F", x"1D", x"1C", x"1A", x"17",
	x"16", x"14", x"11", x"0F", x"0C", x"0A", x"06", x"04", x"00", x"FE", x"FA", x"F8",
	x"F5", x"F1", x"EF", x"EC", x"E8", x"E7", x"E3", x"E2", x"E0", x"DD", x"DC", x"DA",
	x"DA", x"D8", x"D9", x"D8", x"D9", x"D9", x"DB", x"DB", x"DD", x"DF", x"E0", x"E3",
	x"E4", x"E8", x"EB", x"EC", x"F0", x"F3", x"F5", x"F8", x"FA", x"FE", x"00", x"02",
	x"05", x"07", x"0A", x"0B", x"0F", x"10", x"13", x"14", x"17", x"18", x"1B", x"1B",
	x"1D", x"1E", x"1E", x"20", x"1F", x"21", x"20", x"21", x"20", x"21", x"1F", x"20",
	x"1F", x"1D", x"1D", x"1B", x"18", x"17", x"14", x"12", x"0F", x"0D", x"09", x"07",
	x"04", x"FF", x"FD", x"F9", x"F7", x"F3", x"F1", x"ED", x"EC", x"E8", x"E6", x"E3",
	x"E2", x"E1", x"DE", x"DE", x"DC", x"DD", x"DD", x"DC", x"DD", x"DD", x"DD", x"DF",
	x"DE", x"E0", x"E0", x"E3", x"E3", x"E6", x"E7", x"EA", x"EB", x"EE", x"EF", x"F3",
	x"F5", x"F6", x"FA", x"FC", x"FF", x"01", x"05", x"08", x"0A", x"0D", x"0F", x"11",
	x"14", x"16", x"19", x"1A", x"1D", x"1D", x"20", x"21", x"23", x"23", x"24", x"24",
	x"25", x"24", x"24", x"23", x"21", x"20", x"1D", x"1C", x"1A", x"16", x"15", x"11",
	x"10", x"0D", x"0A", x"07", x"03", x"01", x"FD", x"FB", x"F7", x"F6", x"F2", x"F0",
	x"EE", x"EB", x"EA", x"E8", x"E5", x"E4", x"E3", x"E2", x"DF", x"E0", x"DF", x"DD",
	x"DE", x"DD", x"DE", x"DE", x"DF", x"DF", x"E1", x"E2", x"E2", x"E5", x"E5", x"E8",
	x"E9", x"EC", x"EE", x"F0", x"F2", x"F4", x"F7", x"F9", x"FC", x"FE", x"02", x"05",
	x"08", x"0B", x"0C", x"10", x"12", x"15", x"17", x"19", x"1B", x"1C", x"1E", x"1F",
	x"20", x"21", x"22", x"23", x"23", x"23", x"22", x"22", x"21", x"20", x"1E", x"1C",
	x"1B", x"18", x"17", x"14", x"12", x"10", x"0C", x"0A", x"06", x"04", x"00", x"FF",
	x"FB", x"F9", x"F5", x"F4", x"F0", x"EF", x"ED", x"EB", x"E8", x"E7", x"E5", x"E4",
	x"E2", x"E2", x"E0", x"E0", x"DF", x"DF", x"DE", x"DE", x"DD", x"DF", x"DF", x"DF",
	x"E1", x"E1", x"E3", x"E4", x"E5", x"E8", x"E9", x"EC", x"EE", x"F1", x"F4", x"F6",
	x"FA", x"FC", x"00", x"02", x"06", x"08", x"0C", x"0E", x"11", x"13", x"17", x"18",
	x"1B", x"1C", x"1F", x"1F", x"21", x"21", x"23", x"22", x"22", x"21", x"21", x"20",
	x"1E", x"1E", x"1B", x"1B", x"19", x"17", x"16", x"14", x"11", x"10", x"0D", x"0B",
	x"09", x"06", x"04", x"01", x"00", x"FD", x"FB", x"F8", x"F7", x"F3", x"F2", x"F0",
	x"ED", x"EA", x"E9", x"E6", x"E5", x"E2", x"E2", x"E0", x"DF", x"DF", x"DD", x"DE",
	x"DD", x"DD", x"DE", x"DE", x"E0", x"E0", x"E2", x"E3", x"E5", x"E6", x"E9", x"EC",
	x"EE", x"F1", x"F3", x"F6", x"F9", x"FB", x"FF", x"01", x"04", x"07", x"0A", x"0C",
	x"0F", x"10", x"13", x"14", x"17", x"17", x"1A", x"1B", x"1C", x"1E", x"1D", x"1F",
	x"1E", x"1F", x"1E", x"1F", x"1E", x"1E", x"1D", x"1B", x"1B", x"19", x"19", x"17",
	x"16", x"13", x"12", x"0F", x"0E", x"0C", x"08", x"07", x"03", x"02", x"FF", x"FB",
	x"F9", x"F6", x"F4", x"F0", x"EF", x"EB", x"EA", x"E6", x"E4", x"E3", x"E1", x"E0",
	x"DE", x"DE", x"DD", x"DD", x"DD", x"DD", x"DE", x"DF", x"DF", x"E1", x"E3", x"E4",
	x"E7", x"E8", x"EB", x"EC", x"EE", x"F1", x"F3", x"F6", x"F7", x"F9", x"FD", x"FE",
	x"01", x"04", x"06", x"07", x"0A", x"0B", x"0E", x"0F", x"11", x"14", x"14", x"17",
	x"18", x"1A", x"1B", x"1C", x"1D", x"1D", x"1F", x"1E", x"1F", x"1E", x"1D", x"1E",
	x"1C", x"1C", x"1A", x"19", x"17", x"16", x"13", x"12", x"0F", x"0D", x"0A", x"09",
	x"06", x"03", x"01", x"FE", x"FA", x"F9", x"F5", x"F3", x"F0", x"EF", x"ED", x"EB",
	x"E9", x"E7", x"E6", x"E4", x"E4", x"E2", x"E2", x"E0", x"E0", x"E0", x"DF", x"E0",
	x"E0", x"E0", x"E1", x"E3", x"E4", x"E5", x"E6", x"E9", x"EA", x"ED", x"F0", x"F1",
	x"F4", x"F7", x"F8", x"FC", x"FD", x"01", x"03", x"05", x"06", x"0A", x"0A", x"0D",
	x"0E", x"11", x"11", x"14", x"16", x"16", x"19", x"19", x"1B", x"1C", x"1C", x"1E",
	x"1E", x"1F", x"1F", x"20", x"1E", x"1F", x"1D", x"1B", x"1B", x"18", x"17", x"14",
	x"12", x"0F", x"0D", x"0B", x"07", x"06", x"02", x"00", x"FE", x"FA", x"F8", x"F5",
	x"F2", x"F0", x"ED", x"EC", x"E9", x"E8", x"E7", x"E5", x"E5", x"E4", x"E4", x"E2",
	x"E3", x"E2", x"E3", x"E3", x"E2", x"E3", x"E4", x"E4", x"E5", x"E6", x"E6", x"E7",
	x"E9", x"EA", x"EC", x"EE", x"EF", x"F2", x"F4", x"F6", x"F8", x"FA", x"FD", x"FF",
	x"02", x"04", x"08", x"09", x"0D", x"0E", x"11", x"13", x"15", x"18", x"19", x"1A",
	x"1C", x"1C", x"1E", x"1E", x"1E", x"1F", x"1E", x"1F", x"1E", x"1D", x"1D", x"1C",
	x"19", x"19", x"16", x"15", x"13", x"11", x"0E", x"0C", x"0A", x"07", x"05", x"02",
	x"00", x"FE", x"FA", x"F9", x"F6", x"F4", x"F1", x"F0", x"EE", x"EC", x"EB", x"E8",
	x"E7", x"E7", x"E5", x"E5", x"E3", x"E4", x"E3", x"E3", x"E2", x"E3", x"E2", x"E3",
	x"E3", x"E4", x"E5", x"E5", x"E7", x"E7", x"EA", x"EA", x"ED", x"EE", x"F1", x"F3",
	x"F5", x"F8", x"FA", x"FD", x"00", x"03", x"05", x"08", x"0B", x"0E", x"10", x"13",
	x"14", x"17", x"18", x"1A", x"1B", x"1D", x"1C", x"1E", x"1D", x"1D", x"1D", x"1C",
	x"1C", x"1B", x"19", x"19", x"17", x"16", x"16", x"14", x"13", x"12", x"0F", x"0F",
	x"0C", x"0B", x"09", x"06", x"05", x"03", x"00", x"FE", x"FB", x"F9", x"F7", x"F4",
	x"F3", x"EF", x"EE", x"EC", x"E9", x"E8", x"E7", x"E4", x"E4", x"E2", x"E2", x"E1",
	x"E1", x"E0", x"E1", x"E1", x"E2", x"E3", x"E3", x"E5", x"E6", x"E8", x"E9", x"EC",
	x"ED", x"EE", x"F1", x"F2", x"F5", x"F6", x"FA", x"FB", x"FE", x"00", x"03", x"04",
	x"08", x"09", x"0C", x"0E", x"0F", x"12", x"14", x"14", x"17", x"17", x"19", x"19",
	x"1B", x"1C", x"1C", x"1D", x"1D", x"1D", x"1C", x"1B", x"1B", x"1A", x"18", x"17",
	x"14", x"13", x"12", x"10", x"0E", x"0B", x"0A", x"08", x"07", x"05", x"03", x"01",
	x"FF", x"FC", x"FB", x"F7", x"F6", x"F3", x"F2", x"F0", x"EE", x"EC", x"EA", x"E8",
	x"E7", x"E6", x"E4", x"E3", x"E1", x"E1", x"E0", x"E1", x"E0", x"E2", x"E2", x"E3",
	x"E5", x"E6", x"E8", x"EA", x"EC", x"ED", x"F0", x"F2", x"F4", x"F6", x"F9", x"FA",
	x"FD", x"FE", x"01", x"02", x"05", x"07", x"09", x"0A", x"0D", x"0F", x"0F", x"12",
	x"12", x"15", x"15", x"17", x"17", x"19", x"19", x"19", x"1A", x"1A", x"1B", x"1B",
	x"1A", x"1A", x"19", x"19", x"17", x"17", x"15", x"14", x"12", x"11", x"0F", x"0D",
	x"09", x"08", x"06", x"03", x"01", x"FD", x"FC", x"FA", x"F7", x"F5", x"F3", x"F0",
	x"EF", x"EC", x"EC", x"EA", x"E9", x"E7", x"E5", x"E5", x"E3", x"E4", x"E2", x"E3",
	x"E2", x"E3", x"E3", x"E4", x"E4", x"E5", x"E7", x"E9", x"E9", x"EC", x"ED", x"F0",
	x"F1", x"F4", x"F5", x"F7", x"FA", x"FB", x"FE", x"00", x"02", x"04", x"05", x"06",
	x"09", x"09", x"0C", x"0E", x"0F", x"11", x"12", x"13", x"15", x"17", x"17", x"19",
	x"19", x"1A", x"1A", x"1B", x"1B", x"1B", x"1B", x"1B", x"1A", x"18", x"18", x"16",
	x"15", x"12", x"11", x"0E", x"0D", x"0A", x"08", x"05", x"03", x"FF", x"FE", x"FA",
	x"F9", x"F6", x"F4", x"F2", x"F1", x"EF", x"ED", x"EC", x"EB", x"E9", x"E9", x"E8",
	x"E8", x"E7", x"E6", x"E7", x"E5", x"E6", x"E5", x"E7", x"E6", x"E7", x"E7", x"E8",
	x"E9", x"EA", x"EB", x"EC", x"EC", x"EF", x"F0", x"F1", x"F4", x"F5", x"F8", x"FB",
	x"FD", x"FF", x"02", x"04", x"06", x"09", x"0C", x"0E", x"10", x"11", x"12", x"14",
	x"16", x"16", x"18", x"18", x"1A", x"19", x"1B", x"1B", x"1B", x"1B", x"1B", x"1A",
	x"19", x"18", x"17", x"15", x"14", x"12", x"11", x"0F", x"0E", x"0B", x"0B", x"09",
	x"07", x"04", x"02", x"00", x"FD", x"FB", x"F8", x"F7", x"F4", x"F3", x"F0", x"EF",
	x"EE", x"EB", x"EB", x"E9", x"E9", x"E7", x"E7", x"E5", x"E6", x"E5", x"E6", x"E6",
	x"E5", x"E7", x"E7", x"E8", x"E8", x"EA", x"EA", x"EC", x"EC", x"EE", x"F0", x"F0",
	x"F2", x"F3", x"F6", x"F7", x"F9", x"FB", x"FE", x"FF", x"02", x"04", x"07", x"09",
	x"0C", x"0D", x"10", x"11", x"14", x"15", x"16", x"18", x"18", x"19", x"19", x"1A",
	x"19", x"19", x"1A", x"19", x"19", x"17", x"17", x"15", x"15", x"14", x"11", x"11",
	x"0E", x"0E", x"0B", x"0A", x"07", x"06", x"05", x"02", x"01", x"FE", x"FD", x"FB",
	x"F8", x"F7", x"F4", x"F3", x"F1", x"F0", x"ED", x"ED", x"EA", x"EA", x"E9", x"E7",
	x"E7", x"E5", x"E6", x"E5", x"E5", x"E5", x"E6", x"E5", x"E7", x"E6", x"E8", x"E9",
	x"E9", x"EC", x"EC", x"EF", x"F0", x"F3", x"F5", x"F6", x"F9", x"FA", x"FD", x"FF",
	x"01", x"03", x"05", x"08", x"0A", x"0B", x"0E", x"0E", x"11", x"12", x"14", x"14",
	x"16", x"17", x"17", x"18", x"18", x"19", x"18", x"19", x"17", x"18", x"17", x"15",
	x"15", x"13", x"13", x"11", x"10", x"0E", x"0D", x"0B", x"0A", x"07", x"07", x"05",
	x"03", x"02", x"00", x"FF", x"FC", x"FB", x"F8", x"F8", x"F5", x"F4", x"F1", x"F0",
	x"ED", x"EC", x"EA", x"EA", x"E8", x"E6", x"E7", x"E5", x"E6", x"E4", x"E5", x"E4",
	x"E6", x"E5", x"E7", x"E8", x"E9", x"EA", x"EC", x"EE", x"EF", x"F2", x"F3", x"F6",
	x"F7", x"FA", x"FB", x"FD", x"00", x"00", x"03", x"04", x"07", x"07", x"0A", x"0A",
	x"0C", x"0D", x"0F", x"0F", x"11", x"12", x"13", x"15", x"15", x"16", x"16", x"18",
	x"17", x"18", x"17", x"18", x"18", x"16", x"17", x"15", x"15", x"13", x"11", x"10",
	x"0E", x"0D", x"0A", x"09", x"07", x"04", x"02", x"FF", x"FE", x"FB", x"FA", x"F8",
	x"F6", x"F4", x"F3", x"F1", x"EF", x"EE", x"EC", x"EB", x"E9", x"E9", x"E8", x"E8",
	x"E7", x"E7", x"E7", x"E6", x"E7", x"E6", x"E8", x"E8", x"EA", x"EB", x"EC", x"EC",
	x"EF", x"EF", x"F2", x"F2", x"F5", x"F7", x"F8", x"FA", x"FC", x"FE", x"FF", x"00",
	x"03", x"04", x"07", x"07", x"0A", x"0C", x"0D", x"0E", x"10", x"10", x"12", x"12",
	x"14", x"14", x"16", x"15", x"17", x"17", x"17", x"17", x"17", x"16", x"16", x"14",
	x"15", x"13", x"13", x"11", x"10", x"0F", x"0C", x"0C", x"0A", x"07", x"06", x"03",
	x"02", x"00", x"FC", x"FB", x"F8", x"F7", x"F4", x"F3", x"F2", x"EF", x"EF", x"ED",
	x"EB", x"EB", x"E9", x"EA", x"E9", x"E8", x"E9", x"E7", x"E8", x"E8", x"E8", x"E9",
	x"EA", x"EA", x"EB", x"EC", x"EC", x"EE", x"EE", x"F0", x"F1", x"F3", x"F5", x"F6",
	x"F7", x"FA", x"FB", x"FE", x"FE", x"01", x"02", x"05", x"06", x"09", x"09", x"0C",
	x"0D", x"0F", x"10", x"12", x"12", x"14", x"15", x"16", x"16", x"16", x"18", x"17",
	x"18", x"17", x"17", x"16", x"16", x"15", x"14", x"12", x"12", x"0F", x"0E", x"0D",
	x"0A", x"09", x"06", x"05", x"03", x"00", x"00", x"FD", x"FC", x"FA", x"F8", x"F5",
	x"F4", x"F2", x"F1", x"EF", x"EE", x"EC", x"EC", x"EB", x"EA", x"EB", x"E9", x"E9",
	x"EA", x"E9", x"EA", x"EA", x"E9", x"EB", x"EA", x"EB", x"EB", x"ED", x"ED", x"EF",
	x"EF", x"F1", x"F1", x"F4", x"F5", x"F6", x"F8", x"F9", x"FC", x"FE", x"00", x"02",
	x"04", x"05", x"08", x"09", x"0C", x"0C", x"0F", x"10", x"12", x"12", x"15", x"14",
	x"16", x"17", x"16", x"17", x"16", x"17", x"16", x"16", x"14", x"15", x"13", x"13",
	x"12", x"0F", x"0F", x"0D", x"0C", x"0A", x"09", x"07", x"05", x"04", x"02", x"01",
	x"FE", x"FE", x"FB", x"FA", x"F9", x"F6", x"F6", x"F3", x"F2", x"F1", x"EF", x"EF",
	x"ED", x"ED", x"EB", x"EB", x"E9", x"EA", x"E9", x"E8", x"E8", x"E7", x"E9", x"E8",
	x"E9", x"EA", x"EA", x"EC", x"EC", x"EF", x"EF", x"F2", x"F2", x"F5", x"F6", x"F9",
	x"FA", x"FD", x"FF", x"00", x"03", x"04", x"06", x"07", x"0A", x"0A", x"0C", x"0D",
	x"0F", x"10", x"10", x"13", x"13", x"13", x"15", x"14", x"16", x"15", x"16", x"14",
	x"15", x"14", x"13", x"13", x"12", x"10", x"10", x"0E", x"0E", x"0C", x"0B", x"0A",
	x"08", x"07", x"05", x"04", x"02", x"00", x"FE", x"FD", x"FA", x"FA", x"F8", x"F5",
	x"F5", x"F2", x"F2", x"F1", x"EF", x"ED", x"ED", x"EB", x"EB", x"EB", x"EA", x"E9",
	x"E9", x"E8", x"E9", x"E9", x"EA", x"EA", x"EB", x"EB", x"ED", x"ED", x"EF", x"F1",
	x"F1", x"F3", x"F4", x"F7", x"F8", x"FA", x"FB", x"FE", x"FF", x"02", x"03", x"04",
	x"06", x"07", x"09", x"0A", x"0C", x"0C", x"0E", x"0F", x"11", x"11", x"12", x"12",
	x"14", x"13", x"14", x"14", x"14", x"15", x"13", x"14", x"12", x"13", x"11", x"11",
	x"0F", x"0F", x"0D", x"0D", x"0A", x"0A", x"07", x"07", x"04", x"04", x"01", x"00",
	x"FE", x"FD", x"FA", x"FA", x"F7", x"F6", x"F3", x"F3", x"F0", x"F0", x"EE", x"EC",
	x"EC", x"EA", x"EA", x"E9", x"E9", x"E8", x"E9", x"E9", x"E9", x"EA", x"EA", x"EC",
	x"EC", x"EE", x"EE", x"F0", x"F1", x"F2", x"F4", x"F5", x"F7", x"F9", x"F9", x"FC",
	x"FC", x"FF", x"FF", x"02", x"03", x"05", x"06", x"07", x"09", x"0A", x"0C", x"0D",
	x"0D", x"0F", x"0F", x"11", x"12", x"11", x"13", x"12", x"14", x"13", x"14", x"14",
	x"13", x"14", x"12", x"13", x"11", x"11", x"10", x"0E", x"0E", x"0C", x"0A", x"09",
	x"08", x"05", x"05", x"02", x"01", x"FE", x"FD", x"FA", x"F9", x"F8", x"F5", x"F4",
	x"F2", x"F1", x"EF", x"EF", x"ED", x"ED", x"EC", x"EC", x"EB", x"EA", x"EB", x"EA",
	x"EB", x"EA", x"EC", x"EB", x"ED", x"EC", x"EE", x"EE", x"F0", x"F0", x"F2", x"F3",
	x"F5", x"F5", x"F7", x"F7", x"FA", x"FA", x"FD", x"FD", x"00", x"00", x"03", x"03",
	x"05", x"07", x"08", x"0A", x"0A", x"0D", x"0E", x"0F", x"11", x"12", x"12", x"13",
	x"13", x"15", x"14", x"15", x"15", x"14", x"15", x"14", x"12", x"13", x"10", x"10",
	x"0E", x"0E", x"0C", x"0A", x"09", x"06", x"05", x"03", x"02", x"00", x"FE", x"FD",
	x"FB", x"FA", x"F8", x"F7", x"F5", x"F4", x"F2", x"F2", x"F1", x"F0", x"EF", x"EF",
	x"EE", x"ED", x"ED", x"EC", x"EC", x"EB", x"EC", x"EC", x"EC", x"ED", x"ED", x"EC",
	x"EE", x"EE", x"EF", x"EF", x"F2", x"F3", x"F4", x"F5", x"F7", x"F8", x"FA", x"FC",
	x"FD", x"FF", x"00", x"03", x"03", x"06", x"07", x"09", x"09", x"0C", x"0C", x"0E",
	x"0E", x"10", x"10", x"12", x"12", x"13", x"12", x"14", x"13", x"13", x"12", x"13",
	x"12", x"12", x"11", x"11", x"0F", x"0F", x"0E", x"0B", x"0B", x"08", x"08", x"06",
	x"04", x"03", x"01", x"FF", x"FE", x"FC", x"FB", x"F9", x"F9", x"F7", x"F6", x"F4",
	x"F4", x"F2", x"F2", x"F1", x"EF", x"EF", x"EE", x"EE", x"ED", x"EC", x"ED", x"EB",
	x"EC", x"EC", x"EC", x"ED", x"ED", x"ED", x"EE", x"EE", x"F0", x"F0", x"F2", x"F4",
	x"F4", x"F6", x"F7", x"F9", x"FB", x"FB", x"FE", x"FF", x"02", x"02", x"05", x"06",
	x"08", x"09", x"0B", x"0C", x"0E", x"0E", x"10", x"10", x"11", x"11", x"12", x"12",
	x"13", x"12", x"13", x"12", x"12", x"12", x"10", x"11", x"0F", x"0F", x"0E", x"0C",
	x"0C", x"0B", x"0A", x"09", x"07", x"05", x"05", x"02", x"02", x"00", x"FF", x"FD",
	x"FC", x"F9", x"F9", x"F7", x"F5", x"F5", x"F2", x"F2", x"F1", x"EF", x"EF", x"EE",
	x"EE", x"EC", x"ED", x"EC", x"EC", x"EC", x"EB", x"EC", x"EC", x"ED", x"ED", x"EE",
	x"EE", x"F0", x"F0", x"F1", x"F3", x"F4", x"F6", x"F7", x"F9", x"FB", x"FB", x"FE",
	x"FF", x"00", x"03", x"03", x"06", x"07", x"08", x"0A", x"0A", x"0D", x"0E", x"0D",
	x"0F", x"0F", x"10", x"11", x"11", x"10", x"11", x"10", x"11", x"10", x"11", x"0F",
	x"10", x"0E", x"0F", x"0D", x"0D", x"0C", x"0C", x"0A", x"0A", x"09", x"07", x"07",
	x"05", x"03", x"03", x"00", x"00", x"FD", x"FD", x"FA", x"F9", x"F6", x"F6", x"F3",
	x"F3", x"F0", x"F0", x"EE", x"EE", x"EC", x"ED", x"EB", x"EC", x"EB", x"EC", x"EB",
	x"ED", x"ED", x"EE", x"EF", x"EF", x"F0", x"F0", x"F2", x"F2", x"F5", x"F5", x"F6",
	x"F8", x"F8", x"FB", x"FB", x"FD", x"FE", x"00", x"01", x"02", x"02", x"05", x"05",
	x"07", x"08", x"09", x"0B", x"0B", x"0D", x"0D", x"0E", x"10", x"10", x"11", x"12",
	x"11", x"12", x"11", x"12", x"12", x"11", x"11", x"10", x"10", x"0E", x"0E", x"0D",
	x"0C", x"0A", x"09", x"07", x"06", x"05", x"02", x"02", x"00", x"FE", x"FE", x"FB",
	x"FB", x"F8", x"F8", x"F6", x"F5", x"F3", x"F3", x"F2", x"F1", x"F0", x"EF", x"ED",
	x"EE", x"ED", x"ED", x"EC", x"EC", x"ED", x"ED", x"EE", x"ED", x"EF", x"F0", x"F1",
	x"F1", x"F3", x"F4", x"F5", x"F5", x"F7", x"F9", x"F9", x"FB", x"FC", x"FE", x"FE",
	x"00", x"02", x"02", x"04", x"05", x"05", x"07", x"07", x"0A", x"0A", x"0C", x"0D",
	x"0D", x"0F", x"0E", x"10", x"11", x"10", x"12", x"11", x"12", x"12", x"11", x"11",
	x"10", x"10", x"0E", x"0E", x"0C", x"0C", x"0A", x"0A", x"07", x"07", x"04", x"04",
	x"02", x"00", x"FF", x"FD", x"FC", x"FA", x"F9", x"F7", x"F7", x"F6", x"F4", x"F4",
	x"F2", x"F2", x"F2", x"F0", x"F0", x"EF", x"EF", x"EE", x"EF", x"EE", x"EE", x"ED",
	x"EF", x"EE", x"EF", x"EE", x"EF", x"F1", x"F0", x"F2", x"F2", x"F4", x"F4", x"F7",
	x"F7", x"F9", x"FA", x"FC", x"FE", x"FF", x"01", x"02", x"04", x"05", x"06", x"07",
	x"09", x"09", x"0B", x"0B", x"0D", x"0C", x"0E", x"0E", x"10", x"10", x"10", x"11",
	x"11", x"12", x"11", x"11", x"11", x"10", x"10", x"0E", x"0F", x"0D", x"0C", x"0A",
	x"0A", x"07", x"07", x"05", x"04", x"02", x"01", x"00", x"FE", x"FC", x"FB", x"F9",
	x"F9", x"F8", x"F6", x"F6", x"F4", x"F4", x"F3", x"F3", x"F1", x"F2", x"F1", x"F1",
	x"EF", x"F0", x"EF", x"F0", x"F0", x"EF", x"F0", x"EF", x"F0", x"EF", x"F1", x"F1",
	x"F1", x"F2", x"F2", x"F4", x"F4", x"F6", x"F7", x"F9", x"FB", x"FC", x"FD", x"FF",
	x"00", x"03", x"04", x"06", x"06", x"09", x"0A", x"0A", x"0C", x"0C", x"0D", x"0E",
	x"0E", x"0F", x"0F", x"10", x"10", x"0F", x"10", x"0F", x"0F", x"0F", x"0E", x"0E",
	x"0D", x"0D", x"0B", x"0C", x"0A", x"0A", x"08", x"08", x"06", x"06", x"05", x"03",
	x"03", x"00", x"00", x"FE", x"FD", x"FB", x"FB", x"F9", x"F7", x"F6", x"F5", x"F3",
	x"F3", x"F1", x"F1", x"F0", x"F0", x"EF", x"EF", x"EF", x"EE", x"EF", x"EE", x"EF",
	x"EE", x"EF", x"F0", x"F0", x"F1", x"F1", x"F3", x"F4", x"F4", x"F6", x"F6", x"F8",
	x"F9", x"FB", x"FC", x"FC", x"FF", x"00", x"00", x"03", x"03", x"06", x"07", x"07",
	x"09", x"0A", x"0C", x"0C", x"0D", x"0D", x"0F", x"0E", x"0F", x"0E", x"0F", x"0E",
	x"0F", x"0E", x"0F", x"0E", x"0E", x"0E", x"0D", x"0B", x"0C", x"0A", x"0A", x"09",
	x"07", x"08", x"06", x"05", x"03", x"03", x"01", x"01", x"FF", x"FF", x"FD", x"FB",
	x"FA", x"F8", x"F8", x"F5", x"F5", x"F3", x"F3", x"F1", x"F1", x"F0", x"EF", x"EF",
	x"EF", x"EE", x"EF", x"EE", x"EF", x"EE", x"F0", x"EF", x"F1", x"F1", x"F2", x"F2",
	x"F4", x"F5", x"F5", x"F7", x"F8", x"F8", x"FB", x"FB", x"FD", x"FD", x"FF", x"FF",
	x"02", x"02", x"04", x"04", x"06", x"06", x"08", x"08", x"0A", x"0B", x"0B", x"0D",
	x"0D", x"0E", x"0E", x"0F", x"0F", x"10", x"0F", x"0F", x"0E", x"0F", x"0E", x"0D",
	x"0E", x"0C", x"0C", x"0C", x"0A", x"0A", x"08", x"07", x"05", x"05", x"03", x"02",
	x"01", x"00", x"FE", x"FD", x"FC", x"FA", x"FA", x"F7", x"F7", x"F6", x"F4", x"F4",
	x"F2", x"F2", x"F0", x"F1", x"F0", x"EF", x"EF", x"EE", x"EF", x"EF", x"EE", x"F0",
	x"EF", x"F1", x"F0", x"F2", x"F3", x"F4", x"F5", x"F6", x"F6", x"F8", x"F8", x"FB",
	x"FB", x"FD", x"FD", x"FF", x"00", x"00", x"02", x"02", x"04", x"05", x"05", x"07",
	x"08", x"08", x"09", x"09", x"0B", x"0C", x"0C", x"0D", x"0D", x"0F", x"0F", x"0F",
	x"10", x"0F", x"10", x"0F", x"0E", x"0F", x"0D", x"0D", x"0C", x"0A", x"0A", x"08",
	x"08", x"07", x"04", x"04", x"01", x"01", x"FF", x"FE", x"FD", x"FB", x"FA", x"F9",
	x"F8", x"F6", x"F6", x"F5", x"F5", x"F3", x"F4", x"F2", x"F3", x"F2", x"F2", x"F1",
	x"F1", x"F0", x"F1", x"F0", x"F1", x"F0", x"F1", x"F0", x"F1", x"F2", x"F2", x"F4",
	x"F3", x"F5", x"F6", x"F6", x"F8", x"F9", x"FA", x"FC", x"FC", x"FE", x"FE", x"01",
	x"01", x"03", x"03", x"06", x"06", x"08", x"08", x"0A", x"0A", x"0C", x"0B", x"0D",
	x"0D", x"0E", x"0E", x"0F", x"0E", x"0F", x"0F", x"0F", x"0F", x"0F", x"0D", x"0D",
	x"0D", x"0B", x"0B", x"09", x"09", x"07", x"07", x"05", x"04", x"02", x"02", x"01",
	x"FF", x"FE", x"FD", x"FB", x"FB", x"F9", x"F9", x"F8", x"F7", x"F5", x"F5", x"F3",
	x"F4", x"F3", x"F2", x"F2", x"F1", x"F2", x"F2", x"F2", x"F0", x"F1", x"F1", x"F2",
	x"F2", x"F2", x"F1", x"F3", x"F2", x"F4", x"F4", x"F6", x"F5", x"F8", x"F9", x"FA",
	x"FB", x"FB", x"FD", x"FF", x"FF", x"01", x"02", x"04", x"05", x"05", x"08", x"08",
	x"0A", x"0A", x"0B", x"0B", x"0D", x"0D", x"0D", x"0E", x"0D", x"0E", x"0D", x"0E",
	x"0D", x"0D", x"0D", x"0D", x"0B", x"0C", x"0A", x"0B", x"0A", x"08", x"08", x"06",
	x"07", x"05", x"05", x"03", x"01", x"01", x"FF", x"FF", x"FD", x"FD", x"FB", x"FB",
	x"F8", x"F8", x"F7", x"F5", x"F5", x"F4", x"F4", x"F3", x"F2", x"F2", x"F1", x"F1",
	x"F1", x"F1", x"F0", x"F1", x"F0", x"F1", x"F2", x"F2", x"F2", x"F3", x"F3", x"F5",
	x"F4", x"F6", x"F6", x"F7", x"F9", x"F9", x"FC", x"FC", x"FE", x"FF", x"00", x"01",
	x"03", x"03", x"05", x"05", x"07", x"09", x"09", x"0A", x"0A", x"0C", x"0C", x"0D",
	x"0C", x"0E", x"0E", x"0D", x"0E", x"0D", x"0D", x"0C", x"0D", x"0B", x"0B", x"0A",
	x"0A", x"0A", x"08", x"08", x"07", x"07", x"06", x"04", x"04", x"02", x"02", x"00",
	x"00", x"FF", x"FD", x"FD", x"FC", x"FB", x"FA", x"F7", x"F7", x"F5", x"F5", x"F4",
	x"F4", x"F2", x"F2", x"F1", x"F1", x"F1", x"F0", x"F1", x"F0", x"F1", x"F1", x"F2",
	x"F1", x"F3", x"F2", x"F4", x"F4", x"F6", x"F7", x"F7", x"F9", x"F9", x"FB", x"FC",
	x"FC", x"FE", x"FE", x"00", x"00", x"02", x"03", x"03", x"05", x"05", x"07", x"07",
	x"08", x"09", x"09", x"0A", x"0B", x"0B", x"0C", x"0C", x"0C", x"0D", x"0D", x"0C",
	x"0D", x"0C", x"0D", x"0C", x"0C", x"0B", x"0B", x"0A", x"0A", x"08", x"08", x"07",
	x"06", x"05", x"04", x"03", x"02", x"01", x"FF", x"FE", x"FC", x"FC", x"FA", x"F9",
	x"F9", x"F7", x"F7", x"F5", x"F5", x"F4", x"F3", x"F3", x"F1", x"F2", x"F1", x"F2",
	x"F0", x"F1", x"F1", x"F2", x"F1", x"F2", x"F2", x"F4", x"F3", x"F5", x"F5", x"F6",
	x"F6", x"F8", x"F9", x"F9", x"FB", x"FC", x"FC", x"FE", x"FE", x"00", x"00", x"02",
	x"02", x"04", x"05", x"05", x"07", x"06", x"08", x"08", x"0A", x"09", x"0B", x"0C",
	x"0B", x"0D", x"0C", x"0D", x"0C", x"0D", x"0C", x"0D", x"0C", x"0D", x"0B", x"0C",
	x"0A", x"0A", x"08", x"09", x"07", x"06", x"04", x"04", x"02", x"02", x"01", x"FF",
	x"FF", x"FD", x"FB", x"FB", x"FA", x"F8", x"F8", x"F6", x"F7", x"F5", x"F5", x"F4",
	x"F4", x"F4", x"F2", x"F3", x"F2", x"F3", x"F2", x"F3", x"F3", x"F3", x"F2", x"F3",
	x"F3", x"F4", x"F4", x"F5", x"F5", x"F7", x"F6", x"F8", x"F8", x"FA", x"FA", x"FC",
	x"FD", x"FE", x"FE", x"00", x"00", x"02", x"03", x"03", x"05", x"05", x"07", x"08",
	x"07", x"09", x"0A", x"0B", x"0A", x"0C", x"0B", x"0D", x"0C", x"0C", x"0D", x"0D",
	x"0C", x"0D", x"0B", x"0C", x"0A", x"0B", x"09", x"09", x"08", x"08", x"07", x"05",
	x"05", x"04", x"02", x"02", x"01", x"FE", x"FE", x"FC", x"FC", x"FB", x"F9", x"FA",
	x"F8", x"F8", x"F6", x"F6", x"F5", x"F5", x"F4", x"F4", x"F4", x"F2", x"F3", x"F2",
	x"F3", x"F2", x"F3", x"F2", x"F3", x"F3", x"F4", x"F3", x"F5", x"F4", x"F5", x"F6",
	x"F6", x"F8", x"F9", x"FA", x"FB", x"FC", x"FD", x"FD", x"FF", x"FF", x"00", x"02",
	x"02", x"04", x"04", x"06", x"06", x"08", x"08", x"0A", x"0A", x"0B", x"0B", x"0C",
	x"0C", x"0D", x"0D", x"0D", x"0D", x"0C", x"0C", x"0C", x"0A", x"0B", x"09", x"0A",
	x"09", x"07", x"07", x"06", x"06", x"04", x"04", x"02", x"02", x"01", x"FF", x"FF",
	x"FD", x"FD", x"FC", x"FC", x"FB", x"F9", x"F9", x"F8", x"F8", x"F6", x"F7", x"F5",
	x"F5", x"F5", x"F4", x"F3", x"F3", x"F3", x"F2", x"F3", x"F2", x"F3", x"F2", x"F3",
	x"F4", x"F3", x"F5", x"F5", x"F5", x"F7", x"F7", x"F7", x"F9", x"F9", x"FB", x"FB",
	x"FD", x"FE", x"00", x"00", x"02", x"03", x"03", x"05", x"06", x"06", x"07", x"07",
	x"09", x"09", x"09", x"0A", x"0A", x"0B", x"0A", x"0B", x"0C", x"0B", x"0C", x"0A",
	x"0B", x"0B", x"0B", x"09", x"0A", x"08", x"09", x"07", x"08", x"07", x"05", x"05",
	x"04", x"04", x"02", x"02", x"01", x"00", x"FF", x"FD", x"FD", x"FC", x"FA", x"FA",
	x"F8", x"F8", x"F6", x"F6", x"F5", x"F5", x"F4", x"F4", x"F3", x"F4", x"F2", x"F3",
	x"F2", x"F3", x"F2", x"F3", x"F2", x"F4", x"F3", x"F5", x"F4", x"F6", x"F7", x"F6",
	x"F8", x"F8", x"FA", x"FB", x"FC", x"FC", x"FE", x"FE", x"00", x"00", x"02", x"02",
	x"04", x"04", x"06", x"06", x"06", x"08", x"07", x"09", x"09", x"09", x"0A", x"09",
	x"0B", x"0B", x"0A", x"0B", x"0A", x"0B", x"0A", x"0B", x"0A", x"0A", x"09", x"09",
	x"08", x"08", x"08", x"06", x"06", x"04", x"04", x"02", x"03", x"01", x"01", x"FF",
	x"FE", x"FC", x"FC", x"FA", x"FA", x"F8", x"F9", x"F7", x"F7", x"F6", x"F5", x"F5",
	x"F4", x"F4", x"F3", x"F4", x"F3", x"F4", x"F3", x"F4", x"F3", x"F4", x"F3", x"F5",
	x"F4", x"F6", x"F5", x"F7", x"F6", x"F8", x"F8", x"FA", x"F9", x"FB", x"FB", x"FD",
	x"FD", x"FF", x"FF", x"01", x"01", x"02", x"02", x"04", x"04", x"06", x"07", x"07",
	x"08", x"09", x"08", x"0A", x"09", x"0B", x"0A", x"0B", x"0A", x"0B", x"0B", x"0A",
	x"0B", x"0B", x"09", x"0A", x"09", x"09", x"09", x"07", x"07", x"06", x"06", x"04",
	x"04", x"02", x"02", x"00", x"00", x"FE", x"FE", x"FD", x"FB", x"FB", x"FA", x"F8",
	x"F8", x"F6", x"F6", x"F6", x"F5", x"F5", x"F4", x"F4", x"F3", x"F4", x"F3", x"F4",
	x"F3", x"F4", x"F3", x"F5", x"F5", x"F5", x"F6", x"F6", x"F7", x"F8", x"F7", x"F9",
	x"FA", x"F9", x"FB", x"FB", x"FC", x"FD", x"FE", x"FF", x"FF", x"FF", x"01", x"01",
	x"03", x"03", x"05", x"06", x"06", x"07", x"08", x"09", x"09", x"0A", x"0B", x"0B",
	x"0B", x"0C", x"0C", x"0B", x"0C", x"0B", x"0B", x"0A", x"0A", x"0A", x"09", x"09",
	x"08", x"07", x"06", x"05", x"05", x"04", x"03", x"01", x"01", x"FF", x"FF", x"FE",
	x"FD", x"FD", x"FB", x"FB", x"FA", x"FA", x"F9", x"F7", x"F8", x"F6", x"F7", x"F5",
	x"F6", x"F4", x"F5", x"F4", x"F5", x"F3", x"F4", x"F4", x"F4", x"F5", x"F4", x"F5",
	x"F5", x"F6", x"F6", x"F7", x"F8", x"F8", x"F8", x"FA", x"FA", x"FB", x"FB", x"FD",
	x"FD", x"FE", x"00", x"00", x"02", x"03", x"03", x"04", x"05", x"06", x"07", x"08",
	x"07", x"09", x"08", x"0A", x"09", x"0B", x"0B", x"0B", x"0A", x"0B", x"0B", x"0A",
	x"0B", x"09", x"0A", x"09", x"08", x"08", x"07", x"06", x"06", x"05", x"03", x"03",
	x"01", x"02", x"00", x"00", x"FE", x"FE", x"FC", x"FD", x"FB", x"FB", x"FA", x"FA",
	x"F8", x"F9", x"F7", x"F8", x"F6", x"F7", x"F6", x"F6", x"F5", x"F4", x"F5", x"F5",
	x"F3", x"F4", x"F3", x"F5", x"F4", x"F5", x"F4", x"F6", x"F7", x"F7", x"F7", x"F9",
	x"F8", x"FA", x"FB", x"FB", x"FD", x"FD", x"FF", x"00", x"00", x"02", x"02", x"03",
	x"03", x"05", x"05", x"06", x"06", x"08", x"08", x"08", x"09", x"08", x"09", x"09",
	x"0A", x"09", x"0A", x"09", x"0A", x"09", x"0A", x"09", x"09", x"08", x"08", x"07",
	x"07", x"06", x"06", x"05", x"04", x"04", x"02", x"02", x"00", x"00", x"FE", x"FE",
	x"FE", x"FC", x"FC", x"FA", x"FA", x"F9", x"F9", x"F8", x"F8", x"F6", x"F7", x"F6",
	x"F6", x"F5", x"F5", x"F5", x"F4", x"F5", x"F5", x"F4", x"F5", x"F4", x"F5", x"F5",
	x"F5", x"F6", x"F7", x"F6", x"F8", x"F8", x"FA", x"FA", x"FA", x"FC", x"FC", x"FE",
	x"FE", x"00", x"00", x"02", x"02", x"04", x"04", x"05", x"06", x"06", x"07", x"07",
	x"08", x"08", x"09", x"08", x"09", x"08", x"09", x"09", x"08", x"09", x"08", x"09",
	x"08", x"09", x"07", x"08", x"07", x"07", x"07", x"06", x"06", x"04", x"05", x"04",
	x"02", x"03", x"02", x"00", x"00", x"FE", x"FE", x"FC", x"FC", x"FA", x"FA", x"F8",
	x"F9", x"F7", x"F7", x"F6", x"F6", x"F6", x"F5", x"F4", x"F5", x"F5", x"F4", x"F5",
	x"F4", x"F5", x"F5", x"F6", x"F5", x"F7", x"F7", x"F7", x"F8", x"F8", x"F9", x"FA",
	x"FB", x"FA", x"FC", x"FC", x"FD", x"FD", x"FF", x"FF", x"00", x"00", x"02", x"02",
	x"04", x"03", x"05", x"05", x"06", x"06", x"08", x"07", x"09", x"08", x"09", x"09",
	x"0A", x"0A", x"09", x"09", x"0A", x"08", x"09", x"08", x"09", x"08", x"07", x"06",
	x"07", x"05", x"06", x"05", x"03", x"04", x"03", x"01", x"01", x"FF", x"FF", x"FD",
	x"FE", x"FC", x"FC", x"FA", x"FA", x"F8", x"F9", x"F7", x"F7", x"F6", x"F6", x"F6",
	x"F5", x"F4", x"F5", x"F4", x"F5", x"F5", x"F4", x"F6", x"F6", x"F5", x"F7", x"F6",
	x"F8", x"F7", x"F9", x"F8", x"FA", x"FA", x"FA", x"FC", x"FC", x"FC", x"FD", x"FD",
	x"FF", x"FE", x"00", x"00", x"02", x"02", x"02", x"04", x"04", x"05", x"05", x"07",
	x"07", x"08", x"09", x"08", x"0A", x"09", x"0A", x"09", x"0A", x"09", x"0A", x"09",
	x"09", x"09", x"07", x"08", x"06", x"07", x"05", x"05", x"04", x"04", x"02", x"02",
	x"01", x"01", x"FF", x"FF", x"FE", x"FE", x"FD", x"FC", x"FC", x"FA", x"FA", x"F9",
	x"F9", x"F8", x"F8", x"F8", x"F7", x"F7", x"F6", x"F6", x"F6", x"F5", x"F6", x"F6",
	x"F5", x"F6", x"F5", x"F6", x"F6", x"F7", x"F7", x"F8", x"F7", x"F9", x"F9", x"FA",
	x"FA", x"FB", x"FC", x"FC", x"FE", x"FE", x"FF", x"FF", x"01", x"00", x"02", x"03",
	x"02", x"04", x"04", x"05", x"05", x"07", x"06", x"08", x"08", x"08", x"09", x"08",
	x"0A", x"0A", x"09", x"0A", x"09", x"0A", x"08", x"09", x"07", x"08", x"06", x"07",
	x"05", x"05", x"03", x"04", x"02", x"02", x"01", x"00", x"00", x"FE", x"FE", x"FE",
	x"FC", x"FC", x"FC", x"FA", x"FB", x"F9", x"FA", x"F8", x"F9", x"F7", x"F7", x"F8",
	x"F6", x"F7", x"F6", x"F6", x"F5", x"F6", x"F5", x"F6", x"F5", x"F6", x"F5", x"F7",
	x"F6", x"F7", x"F7", x"F8", x"F8", x"FA", x"FA", x"FA", x"FC", x"FC", x"FE", x"FE",
	x"FF", x"01", x"00", x"02", x"02", x"04", x"04", x"05", x"06", x"05", x"07", x"07",
	x"07", x"08", x"08", x"07", x"09", x"08", x"09", x"08", x"09", x"09", x"08", x"08",
	x"07", x"08", x"07", x"07", x"07", x"05", x"06", x"05", x"03", x"04", x"02", x"02",
	x"01", x"01", x"FF", x"00", x"FF", x"FD", x"FD", x"FD", x"FC", x"FB", x"FA", x"FA",
	x"FA", x"F9", x"F7", x"F8", x"F7", x"F7", x"F6", x"F7", x"F5", x"F6", x"F5", x"F6",
	x"F6", x"F5", x"F6", x"F6", x"F6", x"F7", x"F6", x"F8", x"F7", x"F9", x"F8", x"FA",
	x"FA", x"FC", x"FD", x"FD", x"FE", x"FF", x"00", x"00", x"02", x"01", x"03", x"04",
	x"03", x"05", x"05", x"06", x"07", x"06", x"07", x"08", x"07", x"08", x"07", x"08",
	x"08", x"07", x"08", x"07", x"08", x"07", x"08", x"06", x"07", x"07", x"06", x"06",
	x"05", x"05", x"04", x"04", x"03", x"03", x"01", x"01", x"01", x"FF", x"FF", x"FD",
	x"FD", x"FC", x"FC", x"FA", x"FA", x"FA", x"F9", x"F7", x"F8", x"F6", x"F7", x"F6",
	x"F6", x"F5", x"F6", x"F5", x"F6", x"F6", x"F5", x"F7", x"F6", x"F7", x"F7", x"F8",
	x"F8", x"F8", x"F9", x"FA", x"F9", x"FB", x"FC", x"FB", x"FD", x"FE", x"FD", x"FF",
	x"FF", x"01", x"01", x"01", x"03", x"02", x"04", x"04", x"05", x"05", x"05", x"07",
	x"06", x"07", x"07", x"07", x"08", x"07", x"08", x"07", x"08", x"07", x"08", x"07",
	x"08", x"06", x"07", x"06", x"06", x"06", x"04", x"05", x"04", x"03", x"03", x"01",
	x"02", x"01", x"FF", x"00", x"FE", x"FE", x"FC", x"FC", x"FC", x"FA", x"FA", x"F9",
	x"F9", x"F8", x"F8", x"F7", x"F7", x"F7", x"F6", x"F6", x"F5", x"F6", x"F5", x"F6",
	x"F6", x"F7", x"F7", x"F8", x"F8", x"F9", x"F9", x"F9", x"FA", x"F9", x"FA", x"FB",
	x"FB", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"01", x"00", x"02", x"02",
	x"03", x"03", x"05", x"04", x"06", x"05", x"07", x"06", x"08", x"08", x"07", x"09",
	x"08", x"09", x"09", x"08", x"09", x"07", x"08", x"08", x"06", x"07", x"06", x"06",
	x"05", x"03", x"04", x"02", x"02", x"01", x"01", x"FF", x"FF", x"FE", x"FE", x"FC",
	x"FC", x"FC", x"FA", x"FB", x"F9", x"FA", x"F8", x"F9", x"F8", x"F8", x"F7", x"F8",
	x"F7", x"F6", x"F7", x"F7", x"F6", x"F7", x"F6", x"F7", x"F7", x"F8", x"F7", x"F8",
	x"F8", x"F9", x"F9", x"FA", x"FA", x"FB", x"FB", x"FD", x"FD", x"FE", x"FD", x"FF",
	x"FF", x"00", x"01", x"01", x"02", x"03", x"03", x"04", x"05", x"05", x"06", x"06",
	x"07", x"07", x"08", x"08", x"08", x"08", x"07", x"08", x"07", x"08", x"08", x"07",
	x"08", x"06", x"07", x"05", x"06", x"04", x"05", x"03", x"03", x"02", x"02", x"01",
	x"00", x"00", x"FF", x"FF", x"FE", x"FC", x"FD", x"FB", x"FC", x"FA", x"FB", x"F9",
	x"FA", x"F9", x"F9", x"F9", x"F8", x"F7", x"F8", x"F7", x"F8", x"F6", x"F7", x"F7",
	x"F7", x"F7", x"F6", x"F8", x"F7", x"F8", x"F8", x"F9", x"F8", x"FA", x"F9", x"FB",
	x"FB", x"FC", x"FC", x"FE", x"FF", x"FF", x"FF", x"01", x"01", x"02", x"02", x"04",
	x"04", x"04", x"05", x"05", x"06", x"06", x"07", x"06", x"07", x"07", x"08", x"08",
	x"08", x"07", x"08", x"07", x"07", x"06", x"07", x"05", x"05", x"06", x"04", x"04",
	x"04", x"03", x"03", x"03", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FD", x"FE",
	x"FD", x"FC", x"FC", x"FA", x"FB", x"FA", x"F9", x"F9", x"F9", x"F9", x"F8", x"F7",
	x"F8", x"F6", x"F7", x"F6", x"F7", x"F6", x"F7", x"F6", x"F8", x"F7", x"F8", x"F8",
	x"F9", x"F8", x"FA", x"FA", x"FA", x"FC", x"FB", x"FD", x"FD", x"FE", x"FF", x"FF",
	x"00", x"00", x"02", x"02", x"03", x"04", x"04", x"04", x"05", x"05", x"06", x"05",
	x"07", x"07", x"06", x"07", x"07", x"06", x"07", x"06", x"07", x"07", x"06", x"07",
	x"05", x"05", x"06", x"05", x"05", x"04", x"03", x"04", x"02", x"03", x"02", x"02",
	x"00", x"01", x"FF", x"FF", x"FF", x"FD", x"FD", x"FC", x"FC", x"FA", x"FB", x"FA",
	x"F9", x"F9", x"F8", x"F8", x"F7", x"F8", x"F6", x"F7", x"F6", x"F7", x"F7", x"F6",
	x"F7", x"F6", x"F8", x"F7", x"F8", x"F8", x"F9", x"F9", x"FA", x"FA", x"FC", x"FB",
	x"FD", x"FC", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"02", x"02", x"03",
	x"03", x"04", x"04", x"05", x"05", x"06", x"05", x"06", x"07", x"06", x"07", x"06",
	x"07", x"07", x"07", x"07", x"06", x"07", x"06", x"06", x"05", x"06", x"05", x"04",
	x"04", x"03", x"03", x"03", x"01", x"01", x"00", x"00", x"FE", x"FF", x"FD", x"FD",
	x"FC", x"FC", x"FA", x"FB", x"F9", x"FA", x"F8", x"F9", x"F8", x"F8", x"F8", x"F7",
	x"F8", x"F7", x"F8", x"F7", x"F8", x"F7", x"F8", x"F7", x"F9", x"F9", x"F9", x"F9",
	x"FA", x"F9", x"FB", x"FA", x"FC", x"FC", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"02", x"02", x"03", x"03", x"04", x"04", x"05", x"05",
	x"06", x"05", x"07", x"06", x"07", x"07", x"07", x"06", x"07", x"07", x"07", x"07",
	x"06", x"07", x"06", x"06", x"05", x"04", x"04", x"04", x"03", x"02", x"02", x"00",
	x"00", x"00", x"FE", x"FE", x"FD", x"FD", x"FB", x"FC", x"FB", x"FB", x"F9", x"FA",
	x"F9", x"F9", x"F8", x"F9", x"F7", x"F8", x"F7", x"F8", x"F7", x"F8", x"F7", x"F8",
	x"F7", x"F9", x"F9", x"F8", x"F9", x"F9", x"FA", x"F9", x"FB", x"FA", x"FC", x"FB",
	x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"00", x"02", x"02", x"03",
	x"03", x"04", x"04", x"05", x"06", x"05", x"06", x"06", x"07", x"06", x"07", x"07",
	x"07", x"07", x"06", x"07", x"07", x"06", x"06", x"06", x"05", x"05", x"05", x"04",
	x"04", x"03", x"02", x"02", x"00", x"01", x"00", x"FF", x"FF", x"FE", x"FD", x"FD",
	x"FD", x"FB", x"FC", x"FA", x"FB", x"F9", x"FA", x"F9", x"F9", x"F9", x"F8", x"F9",
	x"F8", x"F8", x"F7", x"F8", x"F7", x"F9", x"F8", x"F9", x"F9", x"F8", x"F9", x"F9",
	x"FA", x"F9", x"FB", x"FB", x"FB", x"FC", x"FC", x"FD", x"FD", x"FE", x"FE", x"00",
	x"FF", x"01", x"00", x"02", x"03", x"02", x"04", x"04", x"04", x"05", x"05", x"06",
	x"06", x"06", x"07", x"06", x"07", x"07", x"06", x"07", x"06", x"07", x"06", x"06",
	x"06", x"04", x"05", x"03", x"04", x"03", x"02", x"03", x"01", x"02", x"00", x"00",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FC", x"FC", x"FC", x"FA", x"FB",
	x"F9", x"FA", x"F9", x"F9", x"F8", x"F9", x"F7", x"F8", x"F7", x"F8", x"F7", x"F8",
	x"F8", x"F7", x"F9", x"F8", x"F9", x"F9", x"FA", x"FB", x"FB", x"FC", x"FB", x"FD",
	x"FC", x"FE", x"FD", x"FF", x"00", x"FF", x"01", x"00", x"02", x"01", x"03", x"02",
	x"04", x"04", x"04", x"05", x"04", x"06", x"06", x"06", x"05", x"06", x"05", x"07",
	x"06", x"05", x"06", x"06", x"05", x"06", x"05", x"05", x"04", x"04", x"04", x"03",
	x"03", x"03", x"01", x"02", x"00", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FC", x"FD", x"FB", x"FC", x"FA", x"FB", x"FA", x"FA", x"F9", x"F9", x"F8", x"F8",
	x"F8", x"F7", x"F8", x"F8", x"F8", x"F7", x"F8", x"F7", x"F9", x"F8", x"F9", x"F9",
	x"FA", x"FA", x"FB", x"FB", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"00",
	x"00", x"01", x"01", x"02", x"02", x"03", x"04", x"04", x"04", x"05", x"04", x"05",
	x"05", x"05", x"06", x"05", x"06", x"06", x"05", x"06", x"05", x"06", x"05", x"06",
	x"05", x"06", x"05", x"04", x"05", x"04", x"04", x"03", x"01", x"02", x"01", x"01",
	x"00", x"FF", x"FE", x"FE", x"FD", x"FD", x"FC", x"FB", x"FB", x"FA", x"FB", x"F9",
	x"FA", x"F9", x"F9", x"F8", x"F9", x"F9", x"F8", x"F9", x"F8", x"F9", x"F8", x"F9",
	x"F8", x"F9", x"F8", x"FA", x"F9", x"FA", x"FA", x"FB", x"FA", x"FC", x"FB", x"FD",
	x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"02", x"02", x"03",
	x"03", x"04", x"03", x"05", x"04", x"05", x"04", x"06", x"05", x"06", x"06", x"06",
	x"06", x"06", x"06", x"06", x"06", x"06", x"05", x"05", x"05", x"05", x"04", x"04",
	x"02", x"03", x"01", x"02", x"00", x"01", x"00", x"FE", x"FF", x"FD", x"FE", x"FD",
	x"FC", x"FC", x"FB", x"FA", x"FA", x"FA", x"F9", x"FA", x"F8", x"F8", x"F9", x"F8",
	x"F9", x"F8", x"F9", x"F9", x"F9", x"FA", x"FA", x"FA", x"FA", x"F9", x"FA", x"FA",
	x"FB", x"FB", x"FB", x"FC", x"FB", x"FD", x"FC", x"FE", x"FD", x"FF", x"FE", x"00",
	x"FF", x"01", x"01", x"01", x"03", x"03", x"03", x"04", x"04", x"05", x"05", x"06",
	x"05", x"06", x"05", x"06", x"05", x"06", x"05", x"06", x"06", x"05", x"06", x"04",
	x"04", x"05", x"03", x"04", x"04", x"03", x"03", x"02", x"02", x"00", x"01", x"FF",
	x"00", x"FE", x"FF", x"FD", x"FE", x"FD", x"FC", x"FC", x"FB", x"FB", x"FB", x"FA",
	x"FA", x"F9", x"FA", x"FA", x"F8", x"F9", x"F8", x"F9", x"F9", x"F9", x"F9", x"F9",
	x"FA", x"F9", x"FA", x"FA", x"FA", x"FB", x"FA", x"FB", x"FC", x"FC", x"FD", x"FD",
	x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"02", x"01", x"03", x"02",
	x"04", x"03", x"05", x"04", x"05", x"06", x"05", x"06", x"05", x"06", x"05", x"06",
	x"06", x"06", x"05", x"06", x"04", x"05", x"04", x"04", x"03", x"03", x"02", x"03",
	x"01", x"02", x"00", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FC", x"FD", x"FB", x"FC", x"FC", x"FB", x"FA", x"FA", x"F9", x"FA", x"F8", x"F9",
	x"F9", x"F9", x"F9", x"F9", x"F8", x"F9", x"F8", x"F9", x"FA", x"FA", x"F9", x"FB",
	x"FA", x"FC", x"FB", x"FC", x"FD", x"FC", x"FE", x"FD", x"FF", x"00", x"FF", x"01",
	x"00", x"01", x"01", x"02", x"03", x"02", x"04", x"03", x"04", x"04", x"05", x"04",
	x"05", x"04", x"06", x"05", x"06", x"06", x"05", x"06", x"06", x"04", x"05", x"04",
	x"05", x"03", x"04", x"03", x"03", x"02", x"02", x"02", x"00", x"01", x"FF", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FC", x"FD", x"FB", x"FC", x"FB", x"FB",
	x"FA", x"FA", x"FA", x"FA", x"FA", x"F8", x"F9", x"F8", x"F9", x"F8", x"F9", x"F8",
	x"F9", x"F9", x"FA", x"FA", x"F9", x"FB", x"FA", x"FC", x"FB", x"FD", x"FC", x"FE",
	x"FE", x"FF", x"FF", x"00", x"FF", x"01", x"01", x"01", x"02", x"02", x"02", x"03",
	x"03", x"03", x"04", x"04", x"03", x"05", x"04", x"05", x"04", x"05", x"05", x"04",
	x"05", x"04", x"05", x"04", x"05", x"04", x"05", x"05", x"03", x"04", x"03", x"03",
	x"02", x"02", x"01", x"01", x"00", x"00", x"00", x"FE", x"FF", x"FD", x"FD", x"FD",
	x"FC", x"FC", x"FB", x"FB", x"FB", x"FA", x"FA", x"F9", x"FA", x"F9", x"FA", x"FA",
	x"FA", x"FA", x"F8", x"FA", x"F9", x"FA", x"F9", x"FA", x"FA", x"FB", x"FB", x"FB",
	x"FB", x"FC", x"FB", x"FD", x"FC", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00",
	x"01", x"01", x"02", x"01", x"03", x"02", x"03", x"03", x"04", x"04", x"03", x"05",
	x"04", x"05", x"05", x"05", x"05", x"05", x"04", x"05", x"04", x"05", x"05", x"04",
	x"05", x"03", x"04", x"03", x"03", x"02", x"03", x"01", x"02", x"01", x"00", x"00",
	x"FF", x"FF", x"FD", x"FE", x"FD", x"FC", x"FC", x"FC", x"FA", x"FB", x"FB", x"FA",
	x"FA", x"F9", x"FA", x"F9", x"FA", x"FA", x"F9", x"FA", x"F9", x"FA", x"F9", x"FA",
	x"FA", x"FB", x"FA", x"FB", x"FA", x"FC", x"FB", x"FC", x"FC", x"FC", x"FD", x"FC",
	x"FE", x"FD", x"FF", x"FE", x"00", x"00", x"00", x"01", x"02", x"02", x"02", x"03",
	x"02", x"04", x"04", x"04", x"05", x"04", x"04", x"05", x"04", x"05", x"06", x"04",
	x"05", x"05", x"04", x"05", x"04", x"04", x"03", x"04", x"03", x"03", x"02", x"02",
	x"02", x"01", x"01", x"01", x"FF", x"00", x"FF", x"FE", x"FE", x"FE", x"FD", x"FD",
	x"FC", x"FC", x"FC", x"FB", x"FB", x"FA", x"FB", x"F9", x"FA", x"F9", x"FA", x"F9",
	x"FA", x"F9", x"FA", x"FA", x"FA", x"FA", x"FA", x"FB", x"FA", x"FB", x"FA", x"FC",
	x"FB", x"FB", x"FD", x"FC", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"00",
	x"01", x"01", x"02", x"01", x"03", x"02", x"03", x"03", x"04", x"04", x"05", x"04",
	x"05", x"04", x"05", x"05", x"05", x"04", x"05", x"04", x"05", x"04", x"04", x"03",
	x"04", x"02", x"03", x"02", x"02", x"02", x"02", x"01", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FC", x"FD", x"FC", x"FB", x"FC", x"FA",
	x"FB", x"FA", x"FB", x"F9", x"FA", x"FA", x"F9", x"FA", x"F9", x"FA", x"F9", x"FA",
	x"F9", x"FA", x"FB", x"FB", x"FA", x"FB", x"FB", x"FC", x"FD", x"FC", x"FE", x"FD",
	x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"00", x"01", x"02", x"01", x"03", x"02",
	x"03", x"04", x"03", x"04", x"03", x"05", x"04", x"05", x"05", x"04", x"05", x"04",
	x"05", x"05", x"04", x"05", x"03", x"04", x"03", x"04", x"02", x"03", x"01", x"02",
	x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD",
	x"FD", x"FD", x"FC", x"FC", x"FC", x"FB", x"FB", x"FA", x"FB", x"F9", x"FA", x"F9",
	x"FA", x"F9", x"FA", x"FA", x"FA", x"FA", x"F9", x"FA", x"FA", x"FB", x"FA", x"FC",
	x"FB", x"FC", x"FD", x"FC", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01",
	x"00", x"02", x"01", x"02", x"02", x"03", x"03", x"02", x"04", x"03", x"04", x"03",
	x"04", x"04", x"04", x"05", x"04", x"05", x"04", x"04", x"04", x"04", x"04", x"04",
	x"03", x"04", x"02", x"03", x"02", x"02", x"02", x"01", x"01", x"01", x"00", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FC", x"FC", x"FC", x"FB", x"FB",
	x"FB", x"FA", x"F9", x"FA", x"F9", x"FA", x"F9", x"F9", x"FA", x"FA", x"FA", x"FB",
	x"FA", x"FB", x"FA", x"FB", x"FB", x"FC", x"FB", x"FD", x"FC", x"FD", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"00", x"FF", x"01", x"01", x"02", x"02", x"02", x"02", x"03",
	x"02", x"03", x"03", x"04", x"04", x"03", x"04", x"03", x"05", x"05", x"05", x"05",
	x"05", x"05", x"04", x"03", x"04", x"03", x"04", x"04", x"02", x"03", x"02", x"02",
	x"01", x"01", x"00", x"01", x"FF", x"00", x"FE", x"FF", x"FD", x"FE", x"FD", x"FD",
	x"FB", x"FC", x"FB", x"FB", x"FB", x"FA", x"FB", x"FA", x"FB", x"F9", x"FA", x"F9",
	x"FA", x"F9", x"FB", x"FA", x"FB", x"FA", x"FB", x"FA", x"FB", x"FC", x"FB", x"FC",
	x"FD", x"FC", x"FD", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"00",
	x"01", x"00", x"02", x"01", x"02", x"03", x"02", x"03", x"04", x"03", x"04", x"04",
	x"03", x"05", x"04", x"05", x"05", x"04", x"05", x"04", x"04", x"04", x"03", x"04",
	x"03", x"03", x"02", x"03", x"01", x"02", x"00", x"01", x"00", x"00", x"00", x"FE",
	x"FF", x"FE", x"FE", x"FD", x"FD", x"FC", x"FD", x"FB", x"FC", x"FB", x"FC", x"FB",
	x"FB", x"FA", x"FB", x"FA", x"FB", x"FB", x"FA", x"FB", x"FA", x"FB", x"FA", x"FB",
	x"FA", x"FB", x"FA", x"FC", x"FB", x"FC", x"FB", x"FD", x"FD", x"FC", x"FE", x"FD",
	x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"01", x"00", x"02", x"01", x"02", x"02",
	x"03", x"02", x"04", x"03", x"04", x"03", x"05", x"04", x"05", x"04", x"05", x"04",
	x"05", x"04", x"04", x"04", x"03", x"04", x"02", x"03", x"02", x"02", x"01", x"01",
	x"01", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD",
	x"FD", x"FC", x"FC", x"FB", x"FC", x"FC", x"FA", x"FB", x"FB", x"FA", x"FB", x"FA",
	x"FB", x"FA", x"FB", x"FA", x"FB", x"FA", x"FB", x"FA", x"FB", x"FC", x"FC", x"FC",
	x"FB", x"FD", x"FD", x"FC", x"FE", x"FD", x"FF", x"FE", x"00", x"00", x"FF", x"01",
	x"00", x"02", x"02", x"02", x"03", x"02", x"03", x"03", x"04", x"03", x"04", x"04",
	x"03", x"04", x"03", x"04", x"03", x"04", x"03", x"04", x"03", x"04", x"02", x"03",
	x"02", x"03", x"02", x"01", x"02", x"01", x"01", x"00", x"01", x"FF", x"00", x"00",
	x"FE", x"FF", x"FE", x"FD", x"FE", x"FD", x"FC", x"FD", x"FB", x"FC", x"FC", x"FB",
	x"FB", x"FA", x"FB", x"FA", x"FB", x"FA", x"FB", x"FB", x"FA", x"FB", x"FA", x"FB",
	x"FA", x"FB", x"FB", x"FC", x"FC", x"FB", x"FD", x"FC", x"FD", x"FD", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"02", x"01", x"03", x"02",
	x"03", x"02", x"04", x"04", x"04", x"03", x"04", x"04", x"03", x"04", x"03", x"04",
	x"03", x"04", x"03", x"03", x"02", x"03", x"02", x"03", x"01", x"02", x"02", x"02",
	x"00", x"01", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FD", x"FE", x"FC",
	x"FC", x"FD", x"FC", x"FB", x"FC", x"FA", x"FB", x"FB", x"FB", x"FA", x"FB", x"FA",
	x"FB", x"FB", x"FA", x"FB", x"FA", x"FB", x"FB", x"FC", x"FC", x"FC", x"FC", x"FC",
	x"FD", x"FC", x"FE", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"01",
	x"01", x"01", x"01", x"02", x"01", x"03", x"02", x"03", x"03", x"02", x"04", x"03",
	x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"03", x"04", x"03", x"03",
	x"02", x"03", x"02", x"02", x"01", x"02", x"00", x"01", x"FF", x"00", x"FF", x"FF",
	x"FE", x"FF", x"FD", x"FE", x"FD", x"FD", x"FD", x"FB", x"FB", x"FC", x"FB", x"FB",
	x"FA", x"FB", x"FB", x"FA", x"FB", x"FA", x"FB", x"FA", x"FB", x"FA", x"FB", x"FA",
	x"FC", x"FC", x"FB", x"FC", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"00", x"00", x"00", x"01", x"00", x"02", x"01", x"02", x"01",
	x"03", x"03", x"02", x"03", x"02", x"04", x"03", x"04", x"04", x"03", x"04", x"03",
	x"04", x"03", x"04", x"03", x"04", x"02", x"03", x"02", x"02", x"01", x"02", x"00",
	x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FD", x"FC",
	x"FD", x"FD", x"FB", x"FC", x"FB", x"FC", x"FC", x"FB", x"FC", x"FA", x"FB", x"FA",
	x"FB", x"FA", x"FB", x"FB", x"FB", x"FC", x"FB", x"FC", x"FB", x"FC", x"FC", x"FC",
	x"FD", x"FD", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"00", x"00", x"FF", x"01",
	x"00", x"01", x"01", x"02", x"02", x"03", x"03", x"02", x"03", x"03", x"04", x"03",
	x"04", x"03", x"04", x"03", x"04", x"04", x"03", x"04", x"03", x"03", x"02", x"03",
	x"02", x"01", x"02", x"02", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FD", x"FE", x"FD", x"FC", x"FD", x"FC", x"FC", x"FB", x"FC", x"FB",
	x"FC", x"FC", x"FB", x"FB", x"FA", x"FB", x"FA", x"FB", x"FA", x"FC", x"FB", x"FC",
	x"FB", x"FC", x"FB", x"FB", x"FC", x"FC", x"FD", x"FC", x"FE", x"FD", x"FE", x"FE",
	x"FF", x"FE", x"00", x"00", x"00", x"01", x"01", x"01", x"02", x"01", x"03", x"02",
	x"03", x"02", x"03", x"04", x"04", x"04", x"03", x"04", x"04", x"04", x"04", x"03",
	x"03", x"03", x"03", x"02", x"03", x"01", x"02", x"01", x"02", x"01", x"01", x"00",
	x"01", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FD", x"FE", x"FE", x"FC",
	x"FD", x"FC", x"FC", x"FB", x"FC", x"FB", x"FC", x"FB", x"FB", x"FB", x"FB", x"FB",
	x"FA", x"FB", x"FA", x"FC", x"FB", x"FC", x"FC", x"FB", x"FC", x"FC", x"FD", x"FC",
	x"FD", x"FD", x"FE", x"FE", x"FD", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"01",
	x"00", x"02", x"01", x"02", x"02", x"03", x"02", x"03", x"02", x"03", x"03", x"04",
	x"03", x"04", x"03", x"04", x"02", x"03", x"03", x"03", x"03", x"02", x"03", x"02",
	x"01", x"02", x"01", x"02", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF",
	x"FE", x"FF", x"FD", x"FE", x"FD", x"FD", x"FC", x"FD", x"FC", x"FC", x"FC", x"FC",
	x"FC", x"FB", x"FA", x"FB", x"FA", x"FB", x"FA", x"FB", x"FB", x"FA", x"FC", x"FB",
	x"FC", x"FC", x"FD", x"FC", x"FD", x"FC", x"FE", x"FE", x"FE", x"FE", x"FF", x"FE",
	x"00", x"FF", x"00", x"00", x"00", x"01", x"00", x"01", x"00", x"02", x"01", x"02",
	x"01", x"03", x"03", x"02", x"03", x"02", x"03", x"04", x"03", x"04", x"03", x"04",
	x"03", x"03", x"02", x"03", x"02", x"03", x"01", x"02", x"02", x"01", x"01", x"01",
	x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FC",
	x"FD", x"FD", x"FD", x"FC", x"FC", x"FB", x"FC", x"FC", x"FB", x"FB", x"FA", x"FB",
	x"FB", x"FB", x"FB", x"FC", x"FB", x"FC", x"FB", x"FC", x"FD", x"FD", x"FC", x"FD",
	x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"01",
	x"01", x"00", x"02", x"01", x"02", x"01", x"02", x"02", x"02", x"03", x"03", x"02",
	x"03", x"02", x"04", x"03", x"04", x"03", x"04", x"03", x"02", x"03", x"02", x"03",
	x"02", x"02", x"01", x"02", x"00", x"01", x"FF", x"00", x"FF", x"FF", x"FE", x"FF",
	x"FD", x"FE", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FC", x"FC", x"FC", x"FB",
	x"FC", x"FB", x"FC", x"FC", x"FB", x"FC", x"FB", x"FC", x"FC", x"FC", x"FB", x"FC",
	x"FB", x"FC", x"FD", x"FC", x"FD", x"FC", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"02", x"01", x"02", x"01",
	x"03", x"03", x"02", x"03", x"02", x"03", x"03", x"02", x"03", x"02", x"03", x"02",
	x"03", x"02", x"03", x"03", x"02", x"02", x"01", x"02", x"01", x"01", x"00", x"01",
	x"01", x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FD", x"FC",
	x"FD", x"FC", x"FD", x"FB", x"FC", x"FB", x"FC", x"FB", x"FC", x"FB", x"FB", x"FC",
	x"FB", x"FB", x"FC", x"FB", x"FC", x"FB", x"FC", x"FB", x"FD", x"FD", x"FD", x"FC",
	x"FD", x"FD", x"FE", x"FD", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"01",
	x"00", x"01", x"02", x"01", x"03", x"03", x"02", x"03", x"02", x"03", x"02", x"03",
	x"02", x"03", x"02", x"03", x"02", x"03", x"02", x"03", x"01", x"02", x"02", x"01",
	x"02", x"02", x"01", x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"FE", x"FF",
	x"FF", x"FF", x"FE", x"FD", x"FE", x"FC", x"FD", x"FD", x"FD", x"FC", x"FB", x"FC",
	x"FB", x"FC", x"FB", x"FC", x"FB", x"FC", x"FC", x"FB", x"FC", x"FB", x"FC", x"FC",
	x"FB", x"FD", x"FD", x"FC", x"FD", x"FD", x"FE", x"FD", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"00", x"00", x"FF", x"01", x"00", x"01", x"02", x"01", x"02", x"02", x"03",
	x"02", x"03", x"02", x"03", x"02", x"03", x"03", x"02", x"03", x"02", x"03", x"02",
	x"03", x"02", x"02", x"01", x"02", x"01", x"02", x"01", x"01", x"00", x"00", x"01",
	x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FD", x"FE", x"FD",
	x"FD", x"FD", x"FC", x"FC", x"FB", x"FC", x"FC", x"FB", x"FC", x"FC", x"FC", x"FB",
	x"FC", x"FB", x"FC", x"FC", x"FC", x"FC", x"FC", x"FD", x"FC", x"FD", x"FD", x"FE",
	x"FD", x"FE", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"00", x"01",
	x"00", x"01", x"01", x"01", x"02", x"01", x"02", x"01", x"03", x"02", x"03", x"02",
	x"03", x"03", x"02", x"03", x"02", x"03", x"02", x"03", x"03", x"02", x"02", x"01",
	x"02", x"01", x"01", x"01", x"00", x"01", x"FF", x"00", x"00", x"FF", x"FE", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FC", x"FD", x"FC", x"FC", x"FC",
	x"FB", x"FC", x"FC", x"FC", x"FB", x"FC", x"FB", x"FC", x"FB", x"FC", x"FC", x"FB",
	x"FD", x"FC", x"FD", x"FC", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"01", x"00", x"02", x"01", x"02",
	x"02", x"01", x"02", x"02", x"03", x"02", x"03", x"03", x"02", x"03", x"02", x"03",
	x"03", x"02", x"03", x"02", x"02", x"01", x"02", x"01", x"01", x"01", x"00", x"01",
	x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FC", x"FD",
	x"FC", x"FD", x"FC", x"FD", x"FC", x"FC", x"FB", x"FC", x"FB", x"FC", x"FB", x"FC",
	x"FB", x"FC", x"FB", x"FC", x"FC", x"FD", x"FC", x"FD", x"FD", x"FD", x"FD", x"FE",
	x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"01", x"00",
	x"01", x"00", x"02", x"01", x"02", x"01", x"02", x"02", x"03", x"03", x"02", x"03",
	x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"03", x"01", x"02", x"01", x"02",
	x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FF",
	x"FD", x"FE", x"FD", x"FE", x"FD", x"FC", x"FD", x"FC", x"FD", x"FC", x"FD", x"FC",
	x"FC", x"FC", x"FB", x"FC", x"FB", x"FC", x"FC", x"FB", x"FC", x"FC", x"FD", x"FC",
	x"FD", x"FD", x"FC", x"FD", x"FC", x"FE", x"FD", x"FE", x"FE", x"FE", x"FF", x"FE",
	x"FF", x"FF", x"00", x"FF", x"01", x"01", x"00", x"02", x"01", x"02", x"01", x"02",
	x"03", x"02", x"03", x"02", x"03", x"02", x"03", x"02", x"03", x"02", x"03", x"02",
	x"02", x"01", x"02", x"01", x"02", x"01", x"01", x"00", x"01", x"01", x"01", x"FF",
	x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FC", x"FD", x"FC", x"FD", x"FC", x"FC", x"FC", x"FB", x"FC", x"FB", x"FC", x"FB",
	x"FC", x"FB", x"FC", x"FB", x"FD", x"FC", x"FD", x"FC", x"FD", x"FC", x"FE", x"FD",
	x"FE", x"FD", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"01", x"00",
	x"01", x"01", x"02", x"02", x"02", x"01", x"02", x"01", x"03", x"02", x"03", x"03",
	x"03", x"03", x"02", x"03", x"01", x"02", x"01", x"02", x"01", x"02", x"01", x"02",
	x"00", x"01", x"00", x"01", x"01", x"FF", x"00", x"FF", x"00", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FD", x"FE", x"FD", x"FD", x"FC", x"FD", x"FD", x"FC", x"FC",
	x"FB", x"FC", x"FC", x"FB", x"FC", x"FB", x"FC", x"FB", x"FC", x"FB", x"FD", x"FC",
	x"FD", x"FC", x"FD", x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"01", x"01", x"00", x"01", x"00", x"02", x"01", x"02", x"01",
	x"02", x"02", x"01", x"02", x"01", x"03", x"02", x"03", x"02", x"03", x"01", x"02",
	x"01", x"02", x"01", x"02", x"02", x"01", x"01", x"00", x"01", x"00", x"01", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FC",
	x"FD", x"FC", x"FD", x"FC", x"FD", x"FB", x"FC", x"FB", x"FC", x"FB", x"FC", x"FB",
	x"FC", x"FB", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"00", x"01",
	x"00", x"01", x"00", x"02", x"02", x"01", x"02", x"01", x"02", x"01", x"01", x"03",
	x"02", x"03", x"03", x"02", x"03", x"01", x"02", x"01", x"02", x"01", x"02", x"02",
	x"00", x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FF", x"FE",
	x"FE", x"FD", x"FE", x"FE", x"FC", x"FD", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD",
	x"FD", x"FC", x"FD", x"FD", x"FD", x"FC", x"FD", x"FD", x"FD", x"FD", x"FC", x"FD",
	x"FD", x"FD", x"FD", x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"01", x"00", x"01", x"01", x"02", x"01", x"02",
	x"01", x"02", x"02", x"01", x"03", x"02", x"03", x"02", x"03", x"02", x"02", x"01",
	x"02", x"01", x"02", x"01", x"02", x"00", x"01", x"00", x"01", x"01", x"FF", x"00",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FD",
	x"FC", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD",
	x"FC", x"FD", x"FC", x"FD", x"FC", x"FD", x"FD", x"FD", x"FE", x"FE", x"FD", x"FE",
	x"FD", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"01",
	x"01", x"00", x"02", x"02", x"01", x"02", x"02", x"01", x"02", x"02", x"02", x"03",
	x"02", x"03", x"02", x"02", x"02", x"01", x"02", x"01", x"02", x"02", x"01", x"01",
	x"01", x"01", x"01", x"FF", x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FD", x"FC", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FC", x"FD", x"FD", x"FD", x"FD", x"FC", x"FC", x"FD", x"FC", x"FD",
	x"FD", x"FC", x"FE", x"FD", x"FE", x"FD", x"FE", x"FF", x"FE", x"FF", x"FE", x"00",
	x"FF", x"00", x"00", x"00", x"01", x"00", x"01", x"00", x"02", x"02", x"02", x"02",
	x"02", x"02", x"02", x"02", x"01", x"02", x"01", x"02", x"01", x"02", x"01", x"02",
	x"02", x"02", x"02", x"02", x"00", x"01", x"00", x"01", x"01", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FD",
	x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD", x"FC",
	x"FD", x"FC", x"FD", x"FD", x"FC", x"FD", x"FC", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"00",
	x"01", x"00", x"02", x"01", x"02", x"02", x"01", x"02", x"01", x"02", x"02", x"01",
	x"02", x"02", x"01", x"02", x"01", x"02", x"01", x"02", x"02", x"02", x"00", x"01",
	x"00", x"01", x"01", x"01", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FE", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FC", x"FD", x"FC", x"FD", x"FC", x"FD", x"FC",
	x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FC", x"FD", x"FC", x"FD", x"FC", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"02", x"01", x"02",
	x"01", x"02", x"01", x"02", x"01", x"02", x"01", x"02", x"01", x"02", x"01", x"02",
	x"02", x"02", x"02", x"00", x"01", x"01", x"00", x"01", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FC", x"FD", x"FC", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD",
	x"FC", x"FD", x"FD", x"FC", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"01", x"00", x"01", x"01", x"01", x"02", x"01", x"02", x"01", x"02", x"02", x"02",
	x"01", x"02", x"01", x"01", x"02", x"01", x"02", x"01", x"02", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FC", x"FD", x"FD", x"FC",
	x"FD", x"FC", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD", x"FD",
	x"FD", x"FE", x"FD", x"FE", x"FE", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"01", x"01", x"01", x"00", x"01", x"01", x"02", x"01",
	x"02", x"01", x"02", x"01", x"01", x"02", x"01", x"02", x"01", x"02", x"02", x"01",
	x"02", x"01", x"02", x"00", x"01", x"01", x"01", x"01", x"FF", x"00", x"FF", x"00",
	x"FF", x"FE", x"FF", x"FE", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FC", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FC",
	x"FD", x"FC", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FF", x"FF", x"FE", x"00", x"00", x"FF", x"00", x"00", x"01", x"00", x"01",
	x"00", x"01", x"00", x"02", x"01", x"02", x"01", x"02", x"02", x"02", x"02", x"02",
	x"01", x"02", x"01", x"02", x"01", x"02", x"01", x"02", x"00", x"01", x"00", x"01",
	x"01", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD",
	x"FC", x"FD", x"FD", x"FD", x"FD", x"FC", x"FD", x"FD", x"FD", x"FD", x"FC", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"FF",
	x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"02", x"01", x"02",
	x"02", x"01", x"02", x"01", x"02", x"01", x"02", x"01", x"02", x"01", x"02", x"00",
	x"01", x"01", x"00", x"01", x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FC", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD",
	x"FC", x"FD", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"01",
	x"00", x"01", x"00", x"01", x"01", x"02", x"01", x"02", x"01", x"02", x"01", x"02",
	x"01", x"02", x"01", x"02", x"01", x"02", x"00", x"01", x"01", x"01", x"00", x"01",
	x"00", x"01", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FD", x"FE", x"FE", x"FD", x"FE", x"FC", x"FC", x"FD", x"FC", x"FD", x"FC",
	x"FD", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD", x"FC", x"FE", x"FD", x"FE", x"FE",
	x"FD", x"FE", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"02",
	x"01", x"02", x"01", x"02", x"01", x"02", x"02", x"01", x"02", x"01", x"02", x"02",
	x"02", x"01", x"00", x"01", x"00", x"01", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE",
	x"FD", x"FE", x"FD", x"FD", x"FC", x"FC", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD",
	x"FD", x"FC", x"FD", x"FD", x"FE", x"FD", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"01",
	x"00", x"01", x"00", x"01", x"00", x"02", x"01", x"02", x"01", x"02", x"01", x"02",
	x"01", x"02", x"02", x"02", x"02", x"02", x"00", x"01", x"00", x"01", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FF", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE", x"FD",
	x"FD", x"FC", x"FD", x"FD", x"FD", x"FD", x"FC", x"FD", x"FC", x"FE", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"FE", x"00", x"FF", x"00",
	x"00", x"FF", x"01", x"01", x"01", x"01", x"01", x"00", x"01", x"00", x"02", x"01",
	x"02", x"02", x"01", x"02", x"01", x"02", x"02", x"02", x"01", x"02", x"00", x"01",
	x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FE", x"FD",
	x"FE", x"FE", x"FE", x"FE", x"FD", x"FC", x"FC", x"FD", x"FC", x"FD", x"FC", x"FD",
	x"FC", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE", x"FD", x"FF", x"FE",
	x"FE", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"01", x"00", x"01",
	x"00", x"01", x"00", x"01", x"00", x"02", x"01", x"02", x"01", x"02", x"00", x"01",
	x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"01", x"01", x"01", x"01",
	x"01", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD",
	x"FD", x"FD", x"FC", x"FD", x"FD", x"FD", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD",
	x"FE", x"FD", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"01", x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01",
	x"01", x"02", x"01", x"02", x"01", x"02", x"02", x"02", x"00", x"01", x"00", x"01",
	x"00", x"01", x"00", x"01", x"01", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FD", x"FD", x"FC", x"FD", x"FC", x"FD", x"FC", x"FD", x"FD", x"FD", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"01",
	x"01", x"01", x"00", x"01", x"00", x"01", x"01", x"00", x"02", x"01", x"02", x"02",
	x"02", x"02", x"02", x"01", x"01", x"01", x"01", x"01", x"00", x"01", x"01", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FE", x"FD", x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD",
	x"FE", x"FD", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"01", x"00",
	x"02", x"02", x"01", x"02", x"01", x"02", x"01", x"02", x"02", x"01", x"00", x"01",
	x"00", x"01", x"01", x"00", x"01", x"FF", x"00", x"00", x"00", x"00", x"00", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE",
	x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FD", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"01", x"00",
	x"01", x"00", x"01", x"00", x"01", x"01", x"01", x"00", x"01", x"01", x"00", x"01",
	x"00", x"01", x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"01", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE",
	x"FD", x"FE", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"01", x"00", x"01", x"01", x"01", x"01", x"00", x"01", x"01", x"00",
	x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"01", x"00", x"01", x"00",
	x"01", x"00", x"01", x"00", x"01", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FF", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"01", x"00", x"01",
	x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"01", x"00", x"01",
	x"00", x"00", x"01", x"00", x"01", x"00", x"00", x"01", x"00", x"01", x"01", x"FF",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"FD", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"00", x"00",
	x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"01",
	x"01", x"01", x"01", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"01", x"01", x"00",
	x"01", x"00", x"01", x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"00",
	x"01", x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE",
	x"FE", x"FF", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01",
	x"01", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01",
	x"01", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"01", x"01",
	x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"01", x"01", x"00", x"01",
	x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"00",
	x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"00",
	x"01", x"00", x"01", x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01",
	x"00", x"01", x"00", x"01", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"01", x"01",
	x"01", x"01", x"00", x"01", x"00", x"01", x"01", x"01", x"00", x"01", x"00", x"01",
	x"01", x"00", x"01", x"00", x"01", x"00", x"00", x"01", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"FF", x"00", x"FF", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00",
	x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"01", x"01", x"00", x"01",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"01", x"01",
	x"00", x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00",
	x"01", x"00", x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FF", x"FF",
	x"FE", x"FF", x"FE", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"01", x"01", x"00", x"01", x"00", x"01", x"01", x"00",
	x"01", x"00", x"01", x"01", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"01",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD",
	x"FE", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"01", x"00",
	x"01", x"00", x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"01", x"00",
	x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"01", x"00", x"01", x"01", x"01", x"01", x"00", x"01",
	x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"01", x"00", x"01",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"01",
	x"00", x"01", x"00", x"01", x"00", x"01", x"01", x"01", x"01", x"00", x"01", x"00",
	x"01", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01",
	x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FD", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD",
	x"FE", x"FD", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"01",
	x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01",
	x"01", x"00", x"01", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"01", x"01", x"00", x"01", x"01", x"00", x"01", x"01",
	x"01", x"00", x"01", x"00", x"01", x"01", x"01", x"00", x"01", x"00", x"01", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"01", x"00", x"01", x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"01",
	x"00", x"01", x"01", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FD",
	x"FE", x"FD", x"FE", x"FD", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"01", x"00", x"01", x"00",
	x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"01",
	x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01",
	x"00", x"01", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"FD", x"FE", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FE", x"FF", x"FE", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"01", x"00",
	x"01", x"00", x"01", x"01", x"00", x"01", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FE", x"FF", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FD", x"FE", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"01", x"00", x"01", x"01", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FE", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FD",
	x"FE", x"FD", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"01", x"00", x"01",
	x"01", x"00", x"01", x"00", x"01", x"01", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FD", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FD", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"01", x"01", x"01",
	x"01", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"00", x"01", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"01", x"00", x"01", x"00", x"01", x"01", x"00", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FD", x"FE", x"FD", x"FE", x"FD", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FE", x"FF",
	x"FE", x"FF", x"FF", x"FE", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"01", x"00", x"01", x"01", x"00", x"01",
	x"01", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FD", x"FE",
	x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FD", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"01", x"00", x"01", x"01", x"00", x"01", x"00", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00",
	x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"01", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"00", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FE", x"FF", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FE", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00"
	);
	
signal cnt_out: unsigned(14 downto 0) := (others => '0');	
signal play_sound: std_logic := '0';
constant cnt_max: integer := 15743;
signal out_signal: signed(7 downto 0) := x"00";

begin
	
process (CLK)
begin
    if rising_edge(CLK) then
        if RST = '1' then
            play_sound <= '0';
        elsif PLAY = '1' then
            play_sound <= '1';
        elsif PLAY = '0' and cnt_out = cnt_max then
            play_sound <= '0';
        end if;
    end if;
end process;

	
-- 12bit counter
process (CLK)
begin     
    if rising_edge(CLK) then
        if RST = '1' then
            cnt_out <= (others => '0');
        elsif CE = '1' and play_sound = '1' then
            cnt_out <= cnt_out + 1;       
        end if;
        if cnt_out = cnt_max then
            cnt_out <= (others => '0');            
        end if;        
    end if;
end process;

--SAMPLE_OUT <= kick_sound(conv_integer(cnt_out));
process (CLK) 
begin
    if rising_edge(CLK) then
        if RST = '1' then
            out_signal <= x"00";
        elsif CE = '1' then
            out_signal <= tom2_sound(conv_integer(cnt_out));
        end if;
    end if;    
end process;

SAMPLE_OUT <= out_signal;

end Behavioral;