----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 25.12.2018 17:39:59
-- Design Name: 
-- Module Name: Ride - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Ride is
    Port ( CLK : in STD_LOGIC;
           CE : in STD_LOGIC;
           RST : in STD_LOGIC;
           PLAY : in STD_LOGIC;
           SAMPLE_OUT : out signed(7 downto 0)
           );
end Ride;

architecture Behavioral of Ride is

type memory is array (0 to 107519) of signed(7 downto 0);
constant ride_sound: memory := (
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01",
	x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FD", x"FC", x"FC",
	x"FE", x"FE", x"FC", x"FF", x"FF", x"07", x"04", x"03", x"01", x"FF", x"0A", x"FB",
	x"07", x"02", x"01", x"00", x"F9", x"F9", x"F9", x"01", x"FA", x"01", x"FD", x"01",
	x"FE", x"05", x"FF", x"FA", x"03", x"FE", x"FC", x"01", x"FE", x"FC", x"04", x"FE",
	x"FC", x"FE", x"FE", x"FF", x"04", x"0C", x"02", x"01", x"07", x"01", x"04", x"01",
	x"FD", x"FF", x"FB", x"FC", x"FB", x"FC", x"04", x"FB", x"FF", x"FD", x"F8", x"FE",
	x"03", x"00", x"FD", x"00", x"FF", x"00", x"FA", x"FE", x"FB", x"04", x"02", x"FE",
	x"01", x"05", x"06", x"06", x"0A", x"05", x"02", x"00", x"01", x"00", x"F9", x"FE",
	x"FC", x"FA", x"FE", x"F5", x"FE", x"FE", x"FC", x"FE", x"FA", x"FF", x"FC", x"FD",
	x"00", x"FD", x"00", x"02", x"04", x"06", x"00", x"07", x"07", x"04", x"05", x"FF",
	x"07", x"07", x"00", x"00", x"FD", x"FD", x"FD", x"F9", x"FB", x"F8", x"FB", x"00",
	x"FB", x"FD", x"FC", x"FE", x"FF", x"FF", x"FD", x"FD", x"04", x"00", x"FB", x"FE",
	x"04", x"FF", x"03", x"09", x"FF", x"05", x"03", x"06", x"00", x"00", x"08", x"FE",
	x"05", x"FD", x"F7", x"FD", x"00", x"FF", x"FB", x"FC", x"FF", x"FF", x"FE", x"FD",
	x"F8", x"FD", x"FC", x"FA", x"F8", x"FB", x"01", x"01", x"02", x"01", x"03", x"06",
	x"0B", x"06", x"05", x"09", x"02", x"08", x"02", x"FD", x"04", x"FF", x"01", x"FB",
	x"F9", x"FD", x"F9", x"FF", x"FA", x"FB", x"FD", x"F9", x"FC", x"F8", x"F9", x"FB",
	x"FC", x"00", x"FF", x"FE", x"05", x"05", x"07", x"0A", x"08", x"0B", x"05", x"07",
	x"04", x"FF", x"01", x"01", x"FC", x"F9", x"FC", x"F7", x"FF", x"FE", x"FA", x"FD",
	x"00", x"FE", x"FA", x"FC", x"FE", x"FB", x"FD", x"FB", x"F8", x"FE", x"FD", x"05",
	x"03", x"04", x"04", x"04", x"0A", x"04", x"06", x"09", x"05", x"00", x"FE", x"FD",
	x"FE", x"FC", x"FE", x"FE", x"FB", x"FD", x"FD", x"FF", x"FE", x"01", x"FA", x"01",
	x"FC", x"F7", x"FD", x"F8", x"00", x"F9", x"FE", x"FC", x"FE", x"07", x"04", x"09",
	x"06", x"07", x"08", x"06", x"06", x"00", x"FF", x"05", x"FA", x"F9", x"FE", x"FD",
	x"00", x"FD", x"FB", x"FC", x"FC", x"FD", x"FE", x"FE", x"FD", x"FC", x"FE", x"FD",
	x"FA", x"FB", x"02", x"01", x"01", x"01", x"01", x"07", x"06", x"05", x"03", x"04",
	x"03", x"00", x"03", x"FD", x"FC", x"00", x"FF", x"00", x"FD", x"FE", x"05", x"00",
	x"FD", x"FF", x"FA", x"FD", x"00", x"FA", x"F8", x"FD", x"FD", x"F9", x"FD", x"FF",
	x"00", x"04", x"07", x"FF", x"04", x"08", x"06", x"03", x"03", x"02", x"FD", x"03",
	x"01", x"FC", x"FE", x"05", x"FB", x"FE", x"01", x"FB", x"FF", x"FB", x"FE", x"F9",
	x"F9", x"00", x"FD", x"FE", x"FD", x"FD", x"FF", x"02", x"01", x"FE", x"06", x"07",
	x"01", x"02", x"03", x"FE", x"03", x"04", x"FC", x"FC", x"FF", x"FE", x"FE", x"FD",
	x"00", x"FF", x"03", x"05", x"FB", x"FE", x"03", x"00", x"FB", x"FD", x"FC", x"FF",
	x"00", x"FE", x"FF", x"FE", x"03", x"01", x"00", x"00", x"00", x"FE", x"FF", x"FE",
	x"F9", x"FC", x"02", x"FF", x"FE", x"03", x"00", x"04", x"06", x"04", x"05", x"04",
	x"06", x"02", x"00", x"FD", x"F9", x"FC", x"FC", x"FA", x"F7", x"FC", x"FD", x"FD",
	x"FF", x"FE", x"02", x"02", x"02", x"01", x"FF", x"00", x"FF", x"02", x"00", x"FD",
	x"02", x"00", x"04", x"00", x"01", x"05", x"02", x"03", x"00", x"00", x"01", x"FD",
	x"FD", x"FB", x"FA", x"FB", x"FB", x"02", x"FF", x"FF", x"00", x"00", x"02", x"FF",
	x"01", x"FE", x"00", x"FC", x"FC", x"FC", x"FD", x"00", x"FE", x"02", x"FE", x"01",
	x"05", x"02", x"03", x"08", x"05", x"05", x"02", x"FD", x"00", x"FE", x"FE", x"FA",
	x"F9", x"00", x"FC", x"00", x"FF", x"FE", x"01", x"FD", x"00", x"FA", x"FB", x"FF",
	x"FB", x"FC", x"FA", x"FC", x"02", x"03", x"05", x"04", x"03", x"08", x"08", x"03",
	x"06", x"05", x"01", x"05", x"FE", x"F8", x"FE", x"FD", x"FD", x"FC", x"F9", x"FA",
	x"FA", x"02", x"FB", x"FA", x"FE", x"FE", x"02", x"FA", x"FE", x"FF", x"00", x"04",
	x"FE", x"00", x"04", x"07", x"07", x"04", x"02", x"03", x"04", x"03", x"00", x"FF",
	x"FE", x"01", x"FC", x"FB", x"FC", x"FA", x"03", x"FF", x"FB", x"FD", x"FE", x"FE",
	x"FD", x"FF", x"FA", x"FB", x"00", x"FC", x"FE", x"00", x"FF", x"06", x"06", x"05",
	x"04", x"06", x"08", x"01", x"00", x"00", x"FD", x"FF", x"02", x"FF", x"FD", x"FE",
	x"FF", x"FE", x"FD", x"FF", x"FE", x"00", x"FD", x"FB", x"FC", x"FE", x"FD", x"F9",
	x"FE", x"FD", x"FB", x"FE", x"04", x"02", x"02", x"09", x"04", x"06", x"06", x"03",
	x"03", x"00", x"01", x"FD", x"FF", x"01", x"FC", x"FF", x"FF", x"FE", x"FF", x"00",
	x"00", x"FD", x"FE", x"FE", x"F8", x"F9", x"FA", x"FA", x"FC", x"FE", x"FD", x"FD",
	x"04", x"06", x"04", x"05", x"09", x"09", x"04", x"06", x"FF", x"FE", x"03", x"FD",
	x"FD", x"FA", x"FF", x"FF", x"FE", x"FD", x"FB", x"00", x"03", x"FE", x"FA", x"FD",
	x"FC", x"FD", x"FB", x"FC", x"FB", x"FE", x"03", x"02", x"02", x"02", x"05", x"09",
	x"07", x"04", x"02", x"01", x"03", x"FF", x"F8", x"FA", x"FA", x"FD", x"01", x"FD",
	x"FD", x"00", x"04", x"02", x"FE", x"FE", x"01", x"01", x"FE", x"FA", x"F8", x"FE",
	x"01", x"00", x"FE", x"FE", x"03", x"04", x"04", x"00", x"03", x"05", x"03", x"03",
	x"FC", x"FC", x"FF", x"FD", x"FD", x"FC", x"F9", x"FE", x"04", x"00", x"01", x"03",
	x"01", x"01", x"01", x"FE", x"FD", x"FE", x"FF", x"FC", x"F9", x"FD", x"FF", x"02",
	x"02", x"02", x"02", x"01", x"04", x"FF", x"01", x"01", x"00", x"FE", x"FB", x"FE",
	x"FE", x"FE", x"03", x"01", x"FF", x"04", x"00", x"FF", x"01", x"FF", x"FD", x"FD",
	x"FD", x"FB", x"FE", x"03", x"FE", x"FD", x"01", x"01", x"03", x"02", x"02", x"00",
	x"01", x"00", x"FC", x"FD", x"FF", x"FE", x"FF", x"00", x"FD", x"FE", x"00", x"03",
	x"03", x"00", x"02", x"02", x"FF", x"01", x"FD", x"FA", x"FE", x"FD", x"FC", x"FC",
	x"FD", x"00", x"03", x"06", x"01", x"03", x"08", x"04", x"01", x"FE", x"FD", x"FD",
	x"FE", x"FD", x"FA", x"FB", x"FF", x"FF", x"FE", x"FF", x"FE", x"00", x"05", x"FF",
	x"FF", x"FE", x"00", x"05", x"FE", x"FF", x"00", x"01", x"02", x"03", x"01", x"00",
	x"02", x"03", x"01", x"FE", x"FC", x"FC", x"FF", x"F9", x"F7", x"F9", x"FD", x"01",
	x"FF", x"FE", x"00", x"03", x"05", x"06", x"01", x"03", x"06", x"02", x"01", x"FA",
	x"FE", x"01", x"FF", x"FE", x"FE", x"FE", x"00", x"03", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FC", x"FB", x"FB", x"FE", x"FC", x"FD", x"FF", x"FF", x"05", x"04", x"04",
	x"05", x"02", x"04", x"02", x"00", x"FE", x"FF", x"FD", x"FC", x"FB", x"FB", x"FD",
	x"FE", x"00", x"FF", x"01", x"02", x"03", x"02", x"03", x"03", x"02", x"01", x"FB",
	x"FB", x"FC", x"FC", x"FB", x"FE", x"FF", x"00", x"03", x"FE", x"00", x"01", x"02",
	x"02", x"FF", x"FE", x"FE", x"01", x"FE", x"00", x"01", x"02", x"03", x"03", x"00",
	x"00", x"02", x"FF", x"01", x"FC", x"FA", x"FB", x"FC", x"FD", x"FB", x"FC", x"FD",
	x"FF", x"02", x"02", x"04", x"04", x"04", x"05", x"00", x"FF", x"FF", x"05", x"01",
	x"FD", x"FD", x"FA", x"FD", x"00", x"02", x"FE", x"01", x"04", x"FE", x"FD", x"FE",
	x"FC", x"02", x"FF", x"FC", x"FC", x"FB", x"01", x"00", x"03", x"03", x"01", x"05",
	x"02", x"05", x"FE", x"00", x"02", x"FC", x"FC", x"FA", x"FB", x"FC", x"02", x"FF",
	x"FD", x"01", x"02", x"03", x"02", x"00", x"FF", x"FE", x"01", x"FC", x"FB", x"02",
	x"FF", x"00", x"00", x"FD", x"00", x"02", x"04", x"00", x"02", x"03", x"FE", x"00",
	x"FD", x"FB", x"FE", x"FD", x"FF", x"FB", x"FE", x"00", x"FF", x"00", x"02", x"04",
	x"00", x"03", x"FE", x"FC", x"FF", x"FE", x"FE", x"FE", x"00", x"FF", x"FE", x"03",
	x"03", x"FF", x"06", x"03", x"01", x"00", x"FE", x"00", x"FB", x"00", x"F9", x"FB",
	x"FF", x"FB", x"01", x"FD", x"01", x"02", x"00", x"01", x"FF", x"01", x"03", x"02",
	x"FE", x"FB", x"FF", x"FE", x"FF", x"01", x"00", x"03", x"02", x"03", x"FF", x"00",
	x"05", x"00", x"02", x"FC", x"FA", x"FC", x"FB", x"FE", x"FB", x"FE", x"01", x"FE",
	x"02", x"FE", x"04", x"03", x"01", x"03", x"FC", x"FF", x"FC", x"FD", x"FF", x"FC",
	x"00", x"00", x"04", x"04", x"01", x"05", x"05", x"04", x"01", x"FF", x"FE", x"FD",
	x"00", x"FB", x"FA", x"FC", x"FA", x"FE", x"FB", x"FE", x"FF", x"FF", x"03", x"FD",
	x"00", x"00", x"02", x"03", x"FF", x"03", x"FE", x"FD", x"03", x"00", x"03", x"05",
	x"06", x"04", x"00", x"03", x"FE", x"FE", x"00", x"FC", x"F9", x"F8", x"F8", x"F8",
	x"FD", x"FE", x"FE", x"01", x"02", x"01", x"02", x"03", x"05", x"01", x"03", x"FE",
	x"FC", x"00", x"FF", x"03", x"FF", x"03", x"05", x"FD", x"03", x"04", x"03", x"01",
	x"FF", x"FC", x"F9", x"FD", x"FC", x"FB", x"FD", x"FC", x"FC", x"FD", x"FE", x"01",
	x"04", x"06", x"01", x"01", x"00", x"FE", x"01", x"00", x"00", x"FD", x"00", x"FF",
	x"FD", x"02", x"00", x"04", x"04", x"01", x"02", x"FD", x"01", x"01", x"FE", x"FD",
	x"FB", x"FD", x"FD", x"FE", x"FC", x"FE", x"02", x"02", x"00", x"FF", x"00", x"FF",
	x"00", x"FE", x"F9", x"FB", x"00", x"00", x"00", x"02", x"03", x"05", x"05", x"02",
	x"00", x"06", x"02", x"01", x"00", x"FB", x"FD", x"FB", x"FD", x"FB", x"FC", x"FE",
	x"FF", x"00", x"FD", x"FE", x"00", x"03", x"01", x"FF", x"FE", x"FD", x"FE", x"FE",
	x"FE", x"00", x"03", x"03", x"03", x"02", x"02", x"04", x"05", x"03", x"02", x"FE",
	x"FC", x"00", x"FA", x"F8", x"FE", x"FC", x"FC", x"FE", x"FD", x"00", x"01", x"03",
	x"FF", x"FE", x"00", x"00", x"01", x"00", x"FF", x"00", x"01", x"00", x"00", x"02",
	x"04", x"02", x"01", x"01", x"FD", x"FD", x"FE", x"FE", x"FF", x"FC", x"FB", x"FE",
	x"FC", x"FF", x"02", x"00", x"07", x"04", x"00", x"02", x"01", x"02", x"00", x"01",
	x"FD", x"FC", x"FD", x"F9", x"FB", x"FB", x"FD", x"02", x"00", x"01", x"01", x"03",
	x"04", x"03", x"00", x"00", x"00", x"FD", x"00", x"FE", x"FF", x"03", x"00", x"01",
	x"00", x"00", x"04", x"01", x"00", x"00", x"FB", x"FD", x"FD", x"FD", x"FC", x"FE",
	x"FE", x"FB", x"FF", x"FC", x"01", x"05", x"05", x"04", x"FF", x"00", x"02", x"03",
	x"FF", x"01", x"FF", x"FD", x"00", x"FA", x"FC", x"00", x"03", x"03", x"FD", x"FF",
	x"00", x"01", x"01", x"FE", x"FD", x"FF", x"FF", x"FD", x"FC", x"FF", x"01", x"01",
	x"02", x"FD", x"FF", x"03", x"03", x"01", x"FB", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"01", x"02", x"04", x"00", x"01", x"03", x"04", x"05", x"03", x"FE", x"FA", x"FE",
	x"FE", x"FA", x"FB", x"FD", x"FB", x"FE", x"FC", x"FA", x"00", x"02", x"04", x"00",
	x"02", x"01", x"02", x"03", x"FD", x"FF", x"00", x"02", x"01", x"FE", x"01", x"02",
	x"03", x"03", x"00", x"00", x"01", x"FF", x"FC", x"FA", x"FB", x"FC", x"FC", x"FD",
	x"FF", x"FC", x"00", x"04", x"FF", x"FF", x"02", x"01", x"00", x"00", x"FF", x"FD",
	x"00", x"00", x"FE", x"02", x"00", x"03", x"06", x"02", x"02", x"FF", x"03", x"04",
	x"FF", x"FE", x"FE", x"FD", x"FA", x"FA", x"F9", x"FC", x"FF", x"00", x"FE", x"FC",
	x"00", x"01", x"00", x"01", x"01", x"FF", x"00", x"01", x"FD", x"00", x"03", x"02",
	x"04", x"04", x"01", x"04", x"06", x"02", x"02", x"FE", x"FC", x"FE", x"F9", x"F9",
	x"F9", x"F8", x"FD", x"FD", x"FC", x"FE", x"02", x"06", x"04", x"01", x"00", x"FF",
	x"02", x"00", x"FF", x"FF", x"00", x"02", x"FD", x"00", x"FF", x"03", x"08", x"01",
	x"FF", x"00", x"02", x"FF", x"FF", x"FC", x"FD", x"FF", x"FB", x"FA", x"F9", x"FE",
	x"01", x"02", x"00", x"00", x"00", x"01", x"03", x"00", x"FE", x"FF", x"00", x"FD",
	x"FD", x"FD", x"00", x"04", x"02", x"03", x"00", x"05", x"07", x"03", x"03", x"FE",
	x"FD", x"FD", x"FC", x"F9", x"FA", x"FD", x"FE", x"FC", x"FA", x"FB", x"01", x"04",
	x"02", x"01", x"FF", x"00", x"00", x"00", x"00", x"02", x"04", x"02", x"02", x"FF",
	x"01", x"06", x"03", x"04", x"FE", x"FE", x"FF", x"F9", x"FD", x"F9", x"FB", x"FB",
	x"F8", x"FD", x"FB", x"FF", x"02", x"02", x"03", x"02", x"03", x"05", x"04", x"03",
	x"FE", x"FF", x"FF", x"FC", x"FE", x"FE", x"01", x"00", x"02", x"FF", x"00", x"02",
	x"01", x"03", x"FC", x"FD", x"FC", x"FC", x"FF", x"FA", x"FF", x"01", x"00", x"01",
	x"FD", x"00", x"02", x"01", x"02", x"00", x"00", x"01", x"00", x"FE", x"FC", x"FE",
	x"FE", x"02", x"02", x"FF", x"01", x"03", x"01", x"01", x"02", x"FE", x"FF", x"00",
	x"FB", x"FB", x"FB", x"FD", x"01", x"FE", x"FF", x"FE", x"01", x"05", x"00", x"00",
	x"00", x"01", x"01", x"FC", x"FC", x"FF", x"00", x"00", x"FF", x"FF", x"02", x"06",
	x"07", x"02", x"02", x"FF", x"FD", x"00", x"FB", x"FB", x"FD", x"FD", x"FB", x"F9",
	x"FC", x"FF", x"03", x"03", x"03", x"02", x"00", x"03", x"01", x"01", x"01", x"01",
	x"00", x"FD", x"FE", x"FC", x"00", x"03", x"02", x"FF", x"FF", x"02", x"01", x"01",
	x"00", x"FD", x"FE", x"FF", x"F8", x"FA", x"FD", x"FD", x"00", x"FF", x"00", x"01",
	x"06", x"05", x"04", x"01", x"01", x"00", x"FD", x"FD", x"FE", x"02", x"00", x"00",
	x"FE", x"FD", x"02", x"00", x"02", x"01", x"FE", x"FD", x"FD", x"FD", x"FA", x"FC",
	x"00", x"00", x"FC", x"FF", x"FF", x"00", x"07", x"05", x"05", x"04", x"03", x"01",
	x"FF", x"FF", x"FC", x"FD", x"FF", x"FB", x"F9", x"FC", x"FF", x"01", x"FE", x"00",
	x"02", x"01", x"04", x"00", x"00", x"01", x"00", x"FE", x"FB", x"FF", x"FE", x"00",
	x"02", x"00", x"FE", x"00", x"05", x"00", x"03", x"00", x"FD", x"FE", x"FC", x"FD",
	x"FC", x"FF", x"01", x"FF", x"00", x"FF", x"FD", x"02", x"03", x"02", x"FF", x"FF",
	x"01", x"FD", x"FE", x"FE", x"FE", x"01", x"FF", x"FF", x"FE", x"FF", x"02", x"02",
	x"02", x"00", x"00", x"02", x"02", x"FB", x"FB", x"FE", x"FD", x"FE", x"FE", x"FF",
	x"01", x"01", x"02", x"FF", x"01", x"01", x"00", x"00", x"FE", x"FE", x"FD", x"FE",
	x"00", x"FE", x"FF", x"03", x"01", x"04", x"01", x"01", x"02", x"FF", x"00", x"FD",
	x"FF", x"FF", x"FD", x"FC", x"FA", x"FC", x"FD", x"02", x"00", x"FF", x"02", x"00",
	x"01", x"FF", x"02", x"03", x"02", x"00", x"FC", x"FF", x"FF", x"01", x"02", x"FE",
	x"02", x"03", x"FE", x"01", x"FF", x"00", x"02", x"FF", x"FD", x"F9", x"FD", x"FF",
	x"FD", x"FD", x"FC", x"00", x"00", x"02", x"02", x"02", x"03", x"00", x"00", x"FC",
	x"FF", x"FE", x"01", x"01", x"FE", x"00", x"FF", x"06", x"06", x"02", x"04", x"01",
	x"FE", x"FF", x"FA", x"FB", x"FE", x"FD", x"FB", x"F8", x"FA", x"FA", x"FE", x"01",
	x"FD", x"02", x"03", x"04", x"03", x"02", x"04", x"03", x"03", x"00", x"00", x"00",
	x"01", x"01", x"01", x"02", x"00", x"01", x"00", x"FF", x"FF", x"FB", x"FA", x"FB",
	x"F7", x"FA", x"FB", x"F9", x"FE", x"FE", x"FF", x"01", x"02", x"05", x"06", x"08",
	x"02", x"02", x"04", x"00", x"FF", x"FE", x"00", x"00", x"FF", x"FE", x"FE", x"00",
	x"00", x"01", x"02", x"01", x"FF", x"FF", x"FD", x"FC", x"FC", x"FC", x"FB", x"FD",
	x"FB", x"FC", x"FF", x"FF", x"01", x"01", x"04", x"02", x"02", x"02", x"01", x"02",
	x"FF", x"00", x"00", x"00", x"03", x"02", x"03", x"02", x"01", x"03", x"01", x"01",
	x"FF", x"FD", x"FC", x"F9", x"F6", x"F7", x"FA", x"FA", x"FD", x"FD", x"FD", x"01",
	x"04", x"02", x"02", x"03", x"04", x"05", x"04", x"01", x"01", x"04", x"05", x"02",
	x"FF", x"02", x"04", x"01", x"FF", x"FD", x"FC", x"FF", x"FD", x"FA", x"FA", x"F8",
	x"F8", x"FA", x"F9", x"FB", x"FE", x"02", x"05", x"01", x"03", x"05", x"05", x"06",
	x"04", x"01", x"FF", x"02", x"00", x"FC", x"00", x"FF", x"FF", x"03", x"00", x"00",
	x"01", x"02", x"03", x"FD", x"FB", x"FD", x"FC", x"FD", x"FC", x"F9", x"FB", x"FF",
	x"FF", x"FF", x"03", x"01", x"01", x"00", x"FE", x"FE", x"FF", x"03", x"01", x"01",
	x"01", x"01", x"01", x"02", x"06", x"04", x"04", x"03", x"FF", x"00", x"00", x"FB",
	x"FC", x"FA", x"FA", x"F9", x"F8", x"FC", x"FC", x"FE", x"FE", x"01", x"01", x"01",
	x"05", x"02", x"03", x"01", x"00", x"01", x"00", x"01", x"FE", x"02", x"01", x"00",
	x"03", x"02", x"05", x"03", x"03", x"01", x"FB", x"FB", x"F9", x"FC", x"FC", x"F8",
	x"FB", x"FC", x"FF", x"FF", x"FE", x"02", x"01", x"03", x"03", x"01", x"02", x"FF",
	x"03", x"01", x"FD", x"00", x"FF", x"01", x"FF", x"01", x"FF", x"00", x"05", x"01",
	x"02", x"00", x"FE", x"FE", x"FE", x"FC", x"FA", x"FD", x"00", x"FF", x"FE", x"FC",
	x"FF", x"03", x"01", x"01", x"FF", x"01", x"03", x"FF", x"FE", x"FC", x"FE", x"FF",
	x"01", x"02", x"FE", x"02", x"05", x"02", x"00", x"00", x"03", x"FF", x"00", x"FD",
	x"FA", x"FE", x"FD", x"FD", x"FD", x"00", x"FF", x"01", x"04", x"FF", x"01", x"02",
	x"02", x"03", x"FE", x"FE", x"FF", x"FD", x"FD", x"FA", x"FD", x"FE", x"00", x"01",
	x"FD", x"02", x"FF", x"04", x"05", x"00", x"04", x"01", x"02", x"FE", x"FC", x"00",
	x"FE", x"00", x"FF", x"FF", x"FF", x"01", x"00", x"FE", x"01", x"FE", x"FC", x"FE",
	x"FB", x"FD", x"FE", x"FE", x"FF", x"FF", x"01", x"03", x"03", x"01", x"01", x"02",
	x"00", x"01", x"01", x"00", x"03", x"FF", x"FE", x"FE", x"FF", x"01", x"FF", x"02",
	x"FF", x"FF", x"FE", x"00", x"FF", x"FD", x"FE", x"FD", x"FF", x"FC", x"FB", x"FC",
	x"00", x"01", x"00", x"00", x"01", x"03", x"03", x"02", x"00", x"00", x"FF", x"01",
	x"FF", x"FD", x"01", x"FF", x"02", x"00", x"00", x"03", x"02", x"05", x"00", x"FE",
	x"FD", x"FC", x"FD", x"FC", x"FB", x"FB", x"FB", x"FE", x"FE", x"FD", x"FF", x"03",
	x"04", x"02", x"00", x"00", x"01", x"02", x"01", x"00", x"00", x"01", x"04", x"03",
	x"01", x"FF", x"03", x"04", x"02", x"00", x"FE", x"01", x"FE", x"FB", x"F9", x"F8",
	x"FC", x"FB", x"FB", x"FA", x"FB", x"FE", x"01", x"02", x"02", x"03", x"03", x"05",
	x"02", x"FF", x"00", x"02", x"03", x"01", x"01", x"01", x"04", x"05", x"02", x"01",
	x"01", x"FE", x"00", x"FE", x"F9", x"F9", x"F9", x"F9", x"F8", x"F8", x"FC", x"FF",
	x"FF", x"FF", x"FF", x"02", x"03", x"05", x"04", x"04", x"04", x"04", x"01", x"00",
	x"01", x"01", x"03", x"01", x"00", x"FF", x"03", x"01", x"FD", x"01", x"FF", x"FD",
	x"FC", x"FA", x"F9", x"FB", x"FC", x"FA", x"FD", x"FC", x"00", x"01", x"01", x"03",
	x"02", x"03", x"04", x"03", x"00", x"00", x"01", x"00", x"FE", x"FF", x"FF", x"02",
	x"05", x"02", x"02", x"02", x"02", x"00", x"00", x"FF", x"FC", x"FE", x"FE", x"F9",
	x"F8", x"FB", x"FC", x"FD", x"FD", x"FB", x"FE", x"00", x"00", x"00", x"02", x"04",
	x"05", x"04", x"01", x"01", x"01", x"03", x"04", x"02", x"02", x"02", x"03", x"00",
	x"01", x"FE", x"FC", x"FE", x"FB", x"F8", x"F8", x"FA", x"F9", x"FC", x"FD", x"FB",
	x"FD", x"02", x"05", x"03", x"02", x"03", x"02", x"02", x"02", x"FF", x"02", x"03",
	x"01", x"FF", x"FF", x"02", x"02", x"05", x"02", x"FE", x"FE", x"FD", x"FF", x"FA",
	x"FB", x"FD", x"FC", x"FC", x"FA", x"FC", x"FE", x"02", x"02", x"00", x"03", x"01",
	x"01", x"02", x"00", x"FF", x"FE", x"00", x"00", x"FE", x"00", x"01", x"02", x"02",
	x"01", x"02", x"02", x"04", x"02", x"FE", x"FE", x"FD", x"FD", x"FC", x"FA", x"FB",
	x"FC", x"FE", x"FE", x"FD", x"00", x"04", x"02", x"00", x"00", x"00", x"00", x"FE",
	x"FD", x"FE", x"02", x"02", x"03", x"04", x"02", x"03", x"02", x"02", x"01", x"00",
	x"01", x"FF", x"FA", x"F7", x"FB", x"FA", x"FB", x"FD", x"FB", x"FF", x"02", x"01",
	x"02", x"05", x"06", x"04", x"03", x"00", x"FD", x"FD", x"FF", x"FF", x"FB", x"FD",
	x"FE", x"00", x"03", x"01", x"00", x"03", x"03", x"01", x"FE", x"FF", x"00", x"FE",
	x"FD", x"FA", x"FB", x"FD", x"01", x"02", x"FE", x"02", x"01", x"00", x"00", x"FF",
	x"00", x"01", x"01", x"FC", x"FC", x"FE", x"FE", x"00", x"02", x"01", x"00", x"01",
	x"01", x"02", x"00", x"02", x"00", x"00", x"FE", x"FB", x"FE", x"FD", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"03", x"01", x"01", x"01", x"00", x"03", x"FF", x"FD", x"FE",
	x"FE", x"FF", x"FE", x"FC", x"FE", x"02", x"03", x"00", x"02", x"01", x"FF", x"00",
	x"FC", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"FD", x"04", x"03", x"02", x"03",
	x"01", x"02", x"FD", x"00", x"FE", x"FE", x"00", x"FC", x"FD", x"FA", x"FB", x"FE",
	x"FF", x"00", x"FE", x"01", x"02", x"00", x"01", x"00", x"02", x"03", x"00", x"00",
	x"FF", x"01", x"01", x"00", x"00", x"FE", x"01", x"FE", x"00", x"FF", x"FC", x"00",
	x"FE", x"FB", x"FB", x"FF", x"00", x"FE", x"01", x"FF", x"01", x"04", x"01", x"02",
	x"03", x"02", x"00", x"FE", x"FE", x"FC", x"FC", x"00", x"FF", x"FE", x"FF", x"00",
	x"02", x"01", x"02", x"01", x"03", x"02", x"FF", x"FE", x"FC", x"FF", x"FE", x"FE",
	x"FE", x"FC", x"FF", x"FF", x"FF", x"FD", x"00", x"04", x"01", x"01", x"FD", x"FF",
	x"01", x"FF", x"FF", x"FD", x"FF", x"00", x"00", x"01", x"01", x"04", x"05", x"04",
	x"01", x"FF", x"00", x"FF", x"FD", x"FA", x"F8", x"FB", x"FA", x"FD", x"FE", x"FE",
	x"02", x"FE", x"02", x"00", x"01", x"04", x"02", x"06", x"FF", x"FE", x"FF", x"00",
	x"02", x"00", x"01", x"01", x"01", x"00", x"00", x"01", x"01", x"02", x"FE", x"FA",
	x"FA", x"FA", x"FC", x"FD", x"FC", x"FB", x"FE", x"01", x"00", x"02", x"05", x"03",
	x"04", x"02", x"01", x"02", x"01", x"01", x"FE", x"FE", x"FE", x"FE", x"FF", x"02",
	x"02", x"00", x"02", x"00", x"FE", x"FD", x"FE", x"FE", x"FC", x"FD", x"FA", x"FA",
	x"FE", x"FF", x"00", x"02", x"03", x"01", x"03", x"03", x"00", x"FF", x"05", x"02",
	x"FD", x"00", x"FE", x"00", x"FF", x"FF", x"FF", x"01", x"01", x"FF", x"FE", x"00",
	x"FF", x"FF", x"00", x"FE", x"FB", x"FD", x"FE", x"FC", x"FC", x"FE", x"01", x"01",
	x"02", x"02", x"01", x"04", x"03", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"FD", x"01", x"02", x"FF", x"00", x"03", x"01", x"01", x"FE", x"FA", x"FD", x"FF",
	x"FD", x"FB", x"FC", x"FD", x"FC", x"FF", x"FF", x"FF", x"04", x"04", x"04", x"FE",
	x"FF", x"03", x"02", x"01", x"00", x"01", x"02", x"01", x"00", x"00", x"01", x"02",
	x"01", x"FF", x"FE", x"FD", x"FC", x"FE", x"FB", x"F8", x"FB", x"FB", x"FD", x"FD",
	x"FF", x"00", x"03", x"04", x"02", x"05", x"04", x"04", x"04", x"00", x"FE", x"FD",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"03", x"01", x"FF", x"00", x"00", x"02", x"FF",
	x"FE", x"FB", x"FB", x"FD", x"FA", x"FD", x"FE", x"FF", x"00", x"FF", x"00", x"00",
	x"03", x"06", x"03", x"03", x"01", x"00", x"00", x"FE", x"00", x"FE", x"FF", x"FF",
	x"00", x"01", x"00", x"03", x"02", x"02", x"FF", x"FB", x"FD", x"FE", x"FB", x"FB",
	x"FB", x"FA", x"FD", x"FE", x"00", x"01", x"04", x"03", x"01", x"02", x"01", x"04",
	x"02", x"02", x"FE", x"FC", x"FF", x"FF", x"01", x"00", x"03", x"03", x"01", x"FF",
	x"FD", x"00", x"01", x"FE", x"FD", x"FA", x"FB", x"FB", x"FC", x"FF", x"FD", x"00",
	x"02", x"02", x"02", x"02", x"03", x"04", x"04", x"01", x"FE", x"01", x"FE", x"FF",
	x"FC", x"FC", x"FF", x"FF", x"02", x"FE", x"02", x"02", x"04", x"04", x"FC", x"00",
	x"FF", x"00", x"FE", x"F9", x"FC", x"FD", x"FD", x"FE", x"FF", x"01", x"02", x"03",
	x"00", x"FD", x"FF", x"FF", x"00", x"FF", x"00", x"01", x"01", x"02", x"FF", x"00",
	x"04", x"03", x"01", x"00", x"00", x"FD", x"FE", x"FE", x"FC", x"FE", x"FC", x"FC",
	x"FD", x"FD", x"FE", x"01", x"03", x"03", x"00", x"01", x"02", x"02", x"00", x"00",
	x"FE", x"FE", x"FE", x"FE", x"FD", x"00", x"02", x"00", x"00", x"00", x"02", x"02",
	x"04", x"01", x"FD", x"FF", x"FE", x"FC", x"FD", x"FF", x"FE", x"00", x"01", x"FD",
	x"00", x"02", x"02", x"00", x"00", x"FE", x"FA", x"FE", x"FE", x"FC", x"FF", x"FF",
	x"FF", x"00", x"00", x"02", x"02", x"04", x"05", x"02", x"02", x"00", x"01", x"00",
	x"FE", x"FE", x"FB", x"FF", x"FF", x"FB", x"FC", x"FF", x"00", x"FE", x"FF", x"FD",
	x"FF", x"00", x"FF", x"FD", x"FD", x"00", x"FD", x"01", x"01", x"01", x"04", x"05",
	x"04", x"01", x"02", x"01", x"01", x"00", x"FD", x"FC", x"FB", x"FD", x"FB", x"FE",
	x"FF", x"01", x"02", x"FF", x"00", x"00", x"FF", x"04", x"02", x"FD", x"FF", x"FC",
	x"FE", x"FC", x"FC", x"FE", x"FF", x"01", x"FE", x"FF", x"02", x"03", x"05", x"02",
	x"02", x"FF", x"01", x"02", x"00", x"FF", x"00", x"01", x"FD", x"FF", x"FF", x"02",
	x"02", x"FE", x"FE", x"FD", x"FD", x"FE", x"FB", x"FB", x"FD", x"F9", x"FB", x"FE",
	x"FE", x"01", x"05", x"06", x"04", x"04", x"03", x"04", x"03", x"02", x"01", x"FF",
	x"00", x"FE", x"FD", x"FF", x"00", x"FF", x"FE", x"FF", x"FD", x"FC", x"FF", x"FE",
	x"FB", x"FC", x"FD", x"FE", x"FC", x"FD", x"FE", x"00", x"03", x"01", x"01", x"04",
	x"04", x"04", x"04", x"02", x"01", x"01", x"03", x"FE", x"FE", x"FF", x"FE", x"FF",
	x"FC", x"FF", x"FF", x"01", x"02", x"FF", x"00", x"FD", x"FC", x"FB", x"FB", x"FD",
	x"FA", x"FF", x"00", x"FE", x"FE", x"01", x"03", x"05", x"05", x"02", x"01", x"03",
	x"02", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FC", x"FE", x"01", x"01", x"01",
	x"FE", x"FF", x"FE", x"FD", x"FE", x"FA", x"FD", x"FB", x"FC", x"FD", x"FD", x"01",
	x"00", x"01", x"02", x"03", x"02", x"04", x"05", x"03", x"02", x"00", x"FE", x"FE",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"01", x"02", x"FE", x"FD",
	x"FC", x"FA", x"FD", x"FB", x"FD", x"FE", x"FF", x"00", x"FF", x"01", x"03", x"02",
	x"02", x"02", x"02", x"02", x"FF", x"FF", x"FF", x"01", x"00", x"00", x"01", x"FE",
	x"02", x"01", x"00", x"01", x"FF", x"00", x"FF", x"FC", x"F9", x"FC", x"FC", x"FA",
	x"FD", x"FB", x"FE", x"01", x"02", x"03", x"03", x"04", x"04", x"03", x"02", x"00",
	x"00", x"FF", x"FE", x"FC", x"FB", x"FF", x"01", x"04", x"02", x"FF", x"02", x"00",
	x"00", x"FF", x"FD", x"FE", x"FE", x"FC", x"F9", x"FB", x"FD", x"01", x"03", x"FE",
	x"01", x"01", x"02", x"02", x"00", x"01", x"01", x"00", x"FE", x"FD", x"FF", x"FF",
	x"00", x"01", x"FF", x"00", x"01", x"04", x"02", x"FF", x"00", x"FE", x"FE", x"FD",
	x"FC", x"FE", x"FD", x"FD", x"FF", x"FE", x"00", x"02", x"03", x"04", x"02", x"01",
	x"00", x"01", x"FE", x"FC", x"FD", x"FC", x"FC", x"FD", x"FE", x"00", x"03", x"05",
	x"03", x"04", x"04", x"01", x"FF", x"FF", x"FF", x"FD", x"FD", x"FE", x"FB", x"FE",
	x"FE", x"FE", x"FF", x"00", x"04", x"00", x"01", x"00", x"FF", x"00", x"FE", x"FD",
	x"FC", x"00", x"FE", x"FD", x"00", x"00", x"02", x"03", x"03", x"02", x"02", x"03",
	x"01", x"00", x"00", x"FC", x"FD", x"FE", x"FE", x"FD", x"FE", x"00", x"FD", x"00",
	x"02", x"FF", x"00", x"00", x"01", x"FD", x"FC", x"FE", x"FD", x"01", x"00", x"FF",
	x"FF", x"02", x"03", x"FF", x"02", x"02", x"00", x"02", x"00", x"FC", x"FE", x"FE",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"04", x"02", x"00", x"00", x"02", x"02", x"FD",
	x"FE", x"FB", x"FC", x"FE", x"FD", x"FB", x"FA", x"00", x"01", x"00", x"00", x"01",
	x"04", x"05", x"04", x"01", x"01", x"04", x"01", x"FE", x"FE", x"FC", x"FF", x"00",
	x"FF", x"FF", x"FF", x"02", x"FE", x"FD", x"FC", x"FD", x"FF", x"FC", x"FC", x"FB",
	x"FE", x"FF", x"00", x"03", x"02", x"04", x"01", x"03", x"03", x"00", x"03", x"01",
	x"02", x"FF", x"FD", x"FF", x"FD", x"FF", x"FE", x"FC", x"01", x"FF", x"FF", x"02",
	x"01", x"01", x"FE", x"FF", x"FD", x"FC", x"FF", x"FE", x"FD", x"FC", x"FE", x"00",
	x"02", x"02", x"02", x"04", x"02", x"00", x"FF", x"FF", x"01", x"FF", x"FE", x"FE",
	x"FD", x"FE", x"00", x"03", x"01", x"03", x"05", x"01", x"FF", x"00", x"FE", x"FC",
	x"FC", x"F9", x"FA", x"FB", x"FC", x"FC", x"FD", x"00", x"00", x"03", x"04", x"05",
	x"04", x"02", x"03", x"02", x"01", x"FF", x"00", x"00", x"00", x"FE", x"FC", x"FF",
	x"00", x"00", x"FF", x"FF", x"FE", x"FD", x"FF", x"FC", x"FA", x"FD", x"FD", x"FC",
	x"FE", x"FD", x"01", x"04", x"04", x"04", x"04", x"06", x"05", x"04", x"01", x"FD",
	x"FC", x"FE", x"FE", x"FC", x"FE", x"FE", x"FF", x"00", x"FE", x"FE", x"FF", x"03",
	x"01", x"FF", x"FC", x"FE", x"FF", x"FF", x"FF", x"FC", x"FE", x"01", x"01", x"FF",
	x"00", x"04", x"04", x"05", x"00", x"FE", x"01", x"01", x"FF", x"FD", x"FD", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FA", x"FC", x"FD", x"FE", x"00", x"FF", x"02", x"02", x"03", x"04", x"02", x"04",
	x"03", x"02", x"00", x"FF", x"FD", x"FC", x"FF", x"FE", x"FD", x"FF", x"01", x"FF",
	x"FD", x"FE", x"FE", x"00", x"01", x"FE", x"FE", x"FF", x"FF", x"FD", x"FE", x"01",
	x"01", x"02", x"02", x"00", x"01", x"03", x"04", x"00", x"FF", x"02", x"00", x"FE",
	x"FD", x"FC", x"FD", x"FE", x"FE", x"FD", x"00", x"03", x"01", x"02", x"00", x"FE",
	x"FE", x"00", x"FF", x"FC", x"FD", x"FD", x"FD", x"00", x"FF", x"01", x"04", x"04",
	x"03", x"00", x"02", x"00", x"01", x"02", x"FE", x"FD", x"FD", x"FF", x"FE", x"FC",
	x"FF", x"00", x"02", x"01", x"FF", x"00", x"FF", x"02", x"FD", x"FB", x"FD", x"FC",
	x"FD", x"FE", x"FD", x"FE", x"01", x"05", x"04", x"05", x"05", x"04", x"05", x"02",
	x"01", x"FD", x"FF", x"FE", x"FB", x"FC", x"F9", x"FB", x"FD", x"FF", x"FE", x"FE",
	x"03", x"03", x"02", x"FE", x"FE", x"01", x"FD", x"FE", x"FD", x"FD", x"01", x"04",
	x"02", x"00", x"03", x"05", x"04", x"03", x"FF", x"FE", x"FF", x"FD", x"FC", x"FA",
	x"FE", x"FD", x"FD", x"FE", x"FB", x"00", x"03", x"03", x"02", x"01", x"02", x"FF",
	x"FF", x"FF", x"FD", x"FD", x"FD", x"FF", x"FE", x"FF", x"03", x"04", x"03", x"04",
	x"01", x"01", x"03", x"01", x"FD", x"FC", x"FD", x"FA", x"FC", x"FC", x"FD", x"00",
	x"02", x"01", x"FE", x"02", x"03", x"03", x"02", x"FE", x"FE", x"FD", x"FE", x"FC",
	x"FD", x"01", x"01", x"00", x"00", x"00", x"02", x"03", x"03", x"01", x"FF", x"01",
	x"00", x"FD", x"FC", x"FE", x"FE", x"FE", x"01", x"FC", x"FF", x"02", x"00", x"00",
	x"FF", x"01", x"FE", x"00", x"00", x"FD", x"FF", x"FE", x"00", x"00", x"FF", x"01",
	x"02", x"05", x"02", x"FF", x"01", x"01", x"00", x"FD", x"FD", x"FC", x"FC", x"FE",
	x"FD", x"FD", x"01", x"04", x"04", x"02", x"01", x"FF", x"00", x"00", x"FE", x"FD",
	x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"02", x"04", x"01", x"00", x"00", x"00",
	x"01", x"00", x"FD", x"FD", x"FD", x"FD", x"FD", x"FC", x"FF", x"00", x"01", x"02",
	x"01", x"02", x"04", x"06", x"00", x"FE", x"00", x"FF", x"01", x"FE", x"FD", x"FD",
	x"00", x"FE", x"FD", x"FF", x"01", x"02", x"00", x"00", x"FE", x"FE", x"FF", x"FE",
	x"FD", x"FE", x"FE", x"00", x"01", x"FF", x"02", x"04", x"04", x"03", x"02", x"01",
	x"FF", x"FF", x"FD", x"FD", x"FC", x"FD", x"00", x"FD", x"FE", x"FE", x"01", x"01",
	x"02", x"01", x"00", x"02", x"00", x"FE", x"FD", x"FE", x"FD", x"FE", x"FD", x"FC",
	x"FF", x"02", x"02", x"00", x"04", x"03", x"04", x"04", x"01", x"02", x"00", x"01",
	x"FC", x"FB", x"FE", x"FE", x"00", x"FD", x"FF", x"FF", x"00", x"01", x"FF", x"FF",
	x"FE", x"FD", x"FB", x"FA", x"FD", x"FE", x"00", x"03", x"FF", x"01", x"02", x"04",
	x"05", x"05", x"06", x"03", x"04", x"01", x"FD", x"FF", x"FE", x"FE", x"FC", x"FB",
	x"FB", x"FB", x"FF", x"FE", x"FE", x"FD", x"FD", x"FF", x"FF", x"FE", x"FE", x"00",
	x"00", x"FE", x"00", x"00", x"04", x"04", x"03", x"04", x"02", x"03", x"03", x"04",
	x"01", x"FF", x"FF", x"FB", x"FA", x"FC", x"FC", x"FE", x"00", x"00", x"FF", x"FD",
	x"FF", x"FF", x"00", x"FF", x"FC", x"FD", x"FE", x"FF", x"FD", x"FE", x"01", x"02",
	x"03", x"02", x"03", x"03", x"04", x"04", x"00", x"01", x"02", x"FF", x"FF", x"FE",
	x"FD", x"FD", x"FF", x"FF", x"FB", x"FE", x"00", x"FD", x"FF", x"FD", x"FD", x"FD",
	x"FC", x"FE", x"FC", x"FF", x"FF", x"FF", x"00", x"02", x"04", x"04", x"09", x"06",
	x"04", x"04", x"02", x"FF", x"FF", x"FF", x"FC", x"FD", x"FC", x"FA", x"FB", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FC", x"FF", x"00", x"FE", x"FD",
	x"FE", x"01", x"01", x"04", x"03", x"02", x"03", x"05", x"03", x"00", x"01", x"00",
	x"FF", x"FE", x"FE", x"FD", x"FE", x"00", x"FE", x"FD", x"FF", x"00", x"00", x"01",
	x"FF", x"FD", x"FF", x"FD", x"FA", x"FA", x"FD", x"FC", x"FD", x"01", x"00", x"01",
	x"04", x"06", x"06", x"06", x"06", x"04", x"02", x"01", x"FD", x"FC", x"FF", x"FF",
	x"FD", x"FB", x"FE", x"FD", x"FD", x"00", x"FE", x"00", x"FF", x"FD", x"FB", x"FC",
	x"FF", x"FD", x"FF", x"FF", x"FE", x"00", x"02", x"03", x"04", x"06", x"06", x"04",
	x"03", x"02", x"01", x"01", x"FE", x"FB", x"FB", x"FB", x"FA", x"FC", x"FF", x"FE",
	x"FF", x"FE", x"00", x"01", x"00", x"02", x"01", x"FF", x"FE", x"FE", x"FD", x"FE",
	x"01", x"03", x"02", x"01", x"01", x"02", x"02", x"01", x"00", x"01", x"FE", x"FB",
	x"FB", x"FE", x"FF", x"00", x"00", x"FF", x"00", x"02", x"01", x"01", x"02", x"00",
	x"FF", x"FE", x"FC", x"FE", x"FD", x"FD", x"FE", x"FC", x"FE", x"FF", x"02", x"02",
	x"02", x"04", x"01", x"01", x"02", x"00", x"00", x"FF", x"FF", x"FD", x"FC", x"FC",
	x"FD", x"01", x"00", x"00", x"02", x"01", x"01", x"00", x"FE", x"FE", x"FF", x"FF",
	x"FD", x"FD", x"FC", x"FE", x"02", x"01", x"03", x"02", x"04", x"02", x"FE", x"FF",
	x"FE", x"00", x"FE", x"FD", x"FE", x"FC", x"FF", x"00", x"00", x"00", x"02", x"02",
	x"01", x"01", x"00", x"00", x"00", x"FF", x"FD", x"FD", x"FE", x"FF", x"01", x"FF",
	x"FF", x"00", x"02", x"01", x"01", x"01", x"02", x"FF", x"FD", x"FD", x"FA", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"02", x"01", x"02", x"04", x"04", x"04", x"03", x"FF",
	x"FE", x"FE", x"FF", x"FD", x"FC", x"FD", x"FD", x"00", x"00", x"FF", x"02", x"02",
	x"02", x"FF", x"FF", x"FD", x"FE", x"FF", x"FD", x"FD", x"FD", x"00", x"FE", x"FE",
	x"02", x"01", x"03", x"03", x"03", x"02", x"01", x"03", x"00", x"FF", x"FF", x"FC",
	x"FE", x"00", x"FF", x"FE", x"00", x"01", x"FF", x"FE", x"00", x"FE", x"00", x"00",
	x"FD", x"FA", x"FB", x"FC", x"FE", x"01", x"00", x"02", x"03", x"04", x"02", x"02",
	x"06", x"04", x"02", x"00", x"FE", x"FD", x"FC", x"00", x"FF", x"FE", x"00", x"FE",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FD", x"FB", x"FE", x"FE", x"FD", x"FF",
	x"FC", x"FC", x"00", x"02", x"03", x"04", x"05", x"03", x"04", x"02", x"00", x"02",
	x"03", x"01", x"FC", x"FD", x"FD", x"FD", x"FE", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FD", x"FE", x"01", x"FE", x"FD", x"FB", x"FC", x"FD", x"FF", x"02", x"00", x"05",
	x"05", x"03", x"04", x"02", x"03", x"00", x"02", x"00", x"FD", x"FF", x"FE", x"FE",
	x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"FD", x"FF", x"00", x"FE", x"FC", x"FD",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"02", x"03", x"01", x"00", x"04", x"04", x"04",
	x"03", x"FF", x"00", x"01", x"01", x"FD", x"FD", x"FF", x"FC", x"FE", x"FE", x"FD",
	x"01", x"03", x"00", x"FE", x"FC", x"FD", x"FD", x"FD", x"FE", x"FC", x"FF", x"FF",
	x"00", x"00", x"02", x"05", x"04", x"04", x"02", x"01", x"02", x"03", x"02", x"FE",
	x"00", x"FD", x"FC", x"FF", x"FD", x"FD", x"FE", x"01", x"FF", x"FC", x"00", x"FE",
	x"00", x"FF", x"FB", x"FD", x"FD", x"FF", x"FF", x"FF", x"03", x"00", x"02", x"02",
	x"02", x"03", x"04", x"05", x"01", x"FF", x"FE", x"FC", x"FD", x"FD", x"FE", x"FC",
	x"FE", x"FF", x"FE", x"00", x"00", x"00", x"02", x"01", x"FE", x"FC", x"FE", x"FD",
	x"FE", x"FF", x"FD", x"00", x"00", x"01", x"02", x"02", x"04", x"03", x"02", x"01",
	x"FF", x"01", x"01", x"FF", x"FD", x"FD", x"FF", x"FE", x"FE", x"00", x"00", x"01",
	x"FE", x"FE", x"FE", x"00", x"FF", x"FD", x"FE", x"FC", x"FB", x"FC", x"FF", x"00",
	x"02", x"05", x"04", x"04", x"05", x"04", x"06", x"05", x"01", x"FE", x"FB", x"FC",
	x"FA", x"FA", x"FC", x"FB", x"FF", x"FE", x"FD", x"FE", x"FF", x"03", x"01", x"FF",
	x"FE", x"FF", x"00", x"00", x"00", x"FF", x"00", x"02", x"02", x"01", x"02", x"03",
	x"05", x"02", x"FD", x"FD", x"FF", x"FE", x"FD", x"FC", x"FB", x"FC", x"FD", x"FE",
	x"FD", x"00", x"04", x"02", x"02", x"00", x"00", x"02", x"01", x"00", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FE", x"00", x"01", x"04", x"02", x"01", x"00", x"01", x"00",
	x"FD", x"FD", x"FD", x"FE", x"FF", x"FE", x"FE", x"00", x"02", x"02", x"01", x"01",
	x"00", x"FF", x"00", x"FD", x"FC", x"FC", x"FD", x"FE", x"FD", x"FF", x"01", x"02",
	x"02", x"02", x"02", x"02", x"04", x"03", x"02", x"FF", x"FF", x"FC", x"FD", x"FF",
	x"FC", x"FD", x"FE", x"FD", x"FD", x"FF", x"02", x"01", x"02", x"01", x"FD", x"FE",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"04", x"03", x"FF",
	x"FF", x"FE", x"FE", x"FD", x"FD", x"FE", x"FD", x"FE", x"FF", x"FF", x"00", x"03",
	x"01", x"01", x"02", x"00", x"FF", x"01", x"00", x"FD", x"FC", x"FF", x"FC", x"FD",
	x"01", x"00", x"01", x"03", x"01", x"00", x"01", x"02", x"00", x"01", x"01", x"FC",
	x"FD", x"FE", x"FC", x"FD", x"FE", x"01", x"00", x"00", x"01", x"FF", x"02", x"05",
	x"02", x"FD", x"00", x"FE", x"FC", x"FD", x"FB", x"FF", x"00", x"03", x"00", x"FF",
	x"04", x"03", x"02", x"01", x"FF", x"FE", x"FF", x"FF", x"FB", x"FB", x"FF", x"FE",
	x"FF", x"00", x"FE", x"01", x"02", x"03", x"00", x"FF", x"02", x"01", x"02", x"00",
	x"FF", x"FD", x"FF", x"FE", x"FB", x"00", x"00", x"02", x"01", x"00", x"FE", x"FE",
	x"02", x"FF", x"FD", x"FE", x"FD", x"FE", x"FF", x"FD", x"FF", x"02", x"04", x"03",
	x"01", x"04", x"02", x"03", x"01", x"FE", x"FE", x"FC", x"FD", x"FB", x"FC", x"FC",
	x"FD", x"FF", x"FF", x"01", x"00", x"02", x"02", x"01", x"FF", x"FF", x"00", x"FE",
	x"00", x"FF", x"FE", x"00", x"00", x"00", x"01", x"01", x"03", x"02", x"00", x"00",
	x"FF", x"00", x"FD", x"FE", x"FF", x"FC", x"00", x"FD", x"FD", x"FF", x"FE", x"00",
	x"00", x"02", x"00", x"00", x"00", x"FE", x"FE", x"FF", x"01", x"FF", x"FF", x"FF",
	x"00", x"03", x"02", x"03", x"04", x"02", x"01", x"FE", x"FE", x"FE", x"FD", x"FF",
	x"FD", x"FD", x"FD", x"FD", x"01", x"FE", x"FF", x"FF", x"FD", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"01", x"04", x"03", x"01", x"01", x"02",
	x"03", x"03", x"00", x"FE", x"FF", x"FE", x"FC", x"FB", x"FE", x"FE", x"FE", x"FF",
	x"FC", x"FC", x"01", x"02", x"01", x"FF", x"FE", x"00", x"FF", x"FE", x"FE", x"FD",
	x"01", x"02", x"01", x"01", x"03", x"05", x"04", x"04", x"00", x"FF", x"01", x"00",
	x"FD", x"FB", x"FB", x"FD", x"FE", x"FD", x"FC", x"FE", x"01", x"00", x"FE", x"FE",
	x"FF", x"00", x"01", x"FF", x"FC", x"01", x"00", x"FE", x"00", x"FF", x"01", x"02",
	x"04", x"02", x"01", x"04", x"02", x"02", x"01", x"00", x"FF", x"FE", x"FD", x"FA",
	x"FA", x"FD", x"FC", x"FD", x"01", x"00", x"00", x"00", x"01", x"FE", x"FE", x"00",
	x"FE", x"FE", x"FF", x"FF", x"FE", x"01", x"02", x"01", x"04", x"04", x"02", x"03",
	x"04", x"01", x"00", x"01", x"FE", x"FC", x"FD", x"FD", x"FC", x"FB", x"FC", x"FE",
	x"FF", x"FF", x"FF", x"FE", x"02", x"FE", x"FD", x"FF", x"FF", x"FF", x"FF", x"01",
	x"FE", x"FF", x"03", x"03", x"03", x"04", x"04", x"03", x"04", x"02", x"FE", x"FF",
	x"FF", x"FC", x"FA", x"FB", x"FA", x"F9", x"FD", x"FE", x"FE", x"00", x"02", x"03",
	x"00", x"FF", x"01", x"FF", x"02", x"00", x"FD", x"00", x"00", x"01", x"00", x"01",
	x"01", x"01", x"04", x"00", x"FD", x"00", x"01", x"FF", x"FD", x"FD", x"FD", x"FF",
	x"01", x"FE", x"FE", x"00", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FC",
	x"FB", x"FB", x"00", x"00", x"FE", x"FF", x"00", x"03", x"04", x"03", x"04", x"03",
	x"03", x"00", x"FE", x"FD", x"FD", x"FF", x"FF", x"FE", x"FD", x"01", x"02", x"00",
	x"00", x"FF", x"FF", x"00", x"FD", x"FC", x"FD", x"FD", x"FD", x"FC", x"FD", x"00",
	x"02", x"02", x"02", x"03", x"02", x"04", x"03", x"01", x"01", x"00", x"FF", x"FC",
	x"FD", x"FE", x"FD", x"00", x"FF", x"FF", x"FF", x"01", x"FF", x"FF", x"01", x"FF",
	x"FF", x"00", x"FE", x"FD", x"FD", x"FC", x"FE", x"FE", x"00", x"01", x"03", x"04",
	x"01", x"00", x"01", x"01", x"FF", x"FE", x"FF", x"FC", x"FE", x"00", x"00", x"FF",
	x"03", x"05", x"03", x"02", x"00", x"00", x"FF", x"FF", x"FC", x"F9", x"FD", x"FC",
	x"FA", x"FC", x"FE", x"FE", x"01", x"02", x"01", x"03", x"03", x"03", x"02", x"01",
	x"FF", x"FF", x"01", x"00", x"FD", x"FD", x"FE", x"FF", x"00", x"01", x"01", x"01",
	x"02", x"02", x"FE", x"FE", x"FF", x"00", x"FF", x"FD", x"FB", x"FC", x"FF", x"FF",
	x"FE", x"00", x"02", x"01", x"01", x"01", x"FE", x"00", x"00", x"00", x"FE", x"FE",
	x"FF", x"00", x"02", x"00", x"01", x"04", x"04", x"03", x"01", x"01", x"FF", x"FF",
	x"FE", x"FD", x"FC", x"FC", x"FD", x"FD", x"FD", x"FB", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"02", x"01", x"00", x"00", x"00", x"01", x"02", x"02", x"01", x"03", x"03",
	x"01", x"02", x"02", x"02", x"02", x"01", x"FD", x"FC", x"FC", x"FB", x"FA", x"FB",
	x"FC", x"FD", x"FD", x"FE", x"FF", x"00", x"03", x"02", x"01", x"01", x"00", x"02",
	x"00", x"01", x"00", x"FF", x"02", x"00", x"00", x"00", x"02", x"00", x"01", x"01",
	x"FF", x"01", x"00", x"FF", x"FC", x"FC", x"FC", x"FD", x"00", x"FD", x"FE", x"FF",
	x"FF", x"00", x"FE", x"FE", x"01", x"01", x"00", x"FD", x"FD", x"00", x"FF", x"01",
	x"00", x"01", x"04", x"03", x"05", x"03", x"03", x"03", x"02", x"01", x"FD", x"FE",
	x"FB", x"FC", x"FB", x"FA", x"FC", x"FE", x"00", x"FE", x"FF", x"FF", x"FE", x"01",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"01", x"01", x"04", x"03", x"02",
	x"03", x"02", x"04", x"00", x"FF", x"FF", x"FD", x"FD", x"FD", x"FD", x"FA", x"FD",
	x"FE", x"FD", x"FD", x"00", x"01", x"01", x"01", x"00", x"00", x"01", x"FF", x"FF",
	x"FF", x"FE", x"FD", x"FE", x"01", x"01", x"01", x"05", x"05", x"03", x"01", x"01",
	x"01", x"FF", x"FF", x"FD", x"FC", x"FD", x"FC", x"FD", x"FD", x"FF", x"FF", x"FF",
	x"01", x"FE", x"00", x"02", x"FF", x"FD", x"FE", x"00", x"FE", x"00", x"FF", x"FF",
	x"02", x"02", x"02", x"01", x"04", x"04", x"01", x"02", x"00", x"FE", x"00", x"FF",
	x"FD", x"FD", x"FD", x"FD", x"FC", x"FD", x"FD", x"FF", x"01", x"01", x"00", x"FF",
	x"01", x"FF", x"FD", x"FF", x"FF", x"FE", x"01", x"02", x"FF", x"01", x"04", x"03",
	x"03", x"01", x"01", x"FF", x"00", x"FE", x"FB", x"FD", x"FE", x"FD", x"FD", x"FD",
	x"FE", x"00", x"01", x"01", x"00", x"01", x"02", x"01", x"00", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"01", x"02", x"01", x"FF", x"01", x"01", x"03", x"03", x"01",
	x"00", x"FE", x"FD", x"FC", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"01",
	x"02", x"03", x"01", x"00", x"FF", x"FD", x"FE", x"FD", x"FE", x"FE", x"00", x"00",
	x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"01", x"FF", x"FE", x"FF", x"FE",
	x"00", x"FF", x"00", x"02", x"01", x"02", x"01", x"01", x"00", x"FF", x"FF", x"FE",
	x"FE", x"FD", x"FB", x"FD", x"FD", x"FC", x"FF", x"01", x"01", x"01", x"04", x"03",
	x"01", x"02", x"02", x"01", x"FF", x"FF", x"FC", x"FD", x"FD", x"FA", x"FF", x"01",
	x"02", x"02", x"01", x"03", x"01", x"00", x"00", x"FE", x"FD", x"FD", x"FD", x"FB",
	x"FB", x"00", x"00", x"01", x"00", x"00", x"02", x"02", x"01", x"FF", x"01", x"00",
	x"FD", x"FF", x"FE", x"FF", x"FF", x"01", x"00", x"00", x"03", x"01", x"03", x"02",
	x"FE", x"00", x"FE", x"FE", x"FC", x"FD", x"FF", x"FD", x"FD", x"FC", x"FD", x"00",
	x"00", x"03", x"03", x"01", x"01", x"FF", x"00", x"FE", x"FE", x"00", x"00", x"FF",
	x"FD", x"00", x"02", x"02", x"04", x"02", x"02", x"01", x"01", x"FE", x"FC", x"FE",
	x"FC", x"FC", x"FC", x"FB", x"FE", x"FF", x"00", x"FF", x"01", x"04", x"01", x"03",
	x"01", x"FF", x"00", x"FF", x"FE", x"FD", x"FF", x"FF", x"FF", x"01", x"00", x"FF",
	x"02", x"02", x"02", x"02", x"02", x"00", x"FF", x"FF", x"FB", x"FD", x"FD", x"FF",
	x"FD", x"FC", x"FE", x"FC", x"00", x"01", x"01", x"01", x"00", x"00", x"FC", x"FE",
	x"00", x"00", x"02", x"02", x"01", x"02", x"05", x"03", x"02", x"03", x"02", x"FE",
	x"FE", x"FD", x"FC", x"FC", x"FB", x"FB", x"FA", x"FD", x"FC", x"FF", x"01", x"00",
	x"00", x"00", x"03", x"01", x"02", x"03", x"02", x"01", x"FF", x"00", x"FF", x"01",
	x"02", x"02", x"02", x"00", x"FF", x"00", x"01", x"FE", x"FE", x"FE", x"FD", x"FB",
	x"FA", x"FC", x"FC", x"FF", x"FF", x"00", x"01", x"03", x"02", x"02", x"02", x"00",
	x"01", x"00", x"FF", x"FD", x"FE", x"00", x"00", x"00", x"00", x"03", x"02", x"01",
	x"02", x"00", x"FF", x"FF", x"FF", x"FE", x"FC", x"FC", x"FE", x"FE", x"FE", x"FD",
	x"FE", x"00", x"00", x"00", x"FF", x"00", x"00", x"FE", x"FF", x"FF", x"01", x"01",
	x"03", x"00", x"FE", x"02", x"03", x"03", x"03", x"03", x"02", x"02", x"00", x"FB",
	x"FD", x"FE", x"FC", x"FA", x"FA", x"FA", x"FA", x"FE", x"01", x"00", x"02", x"03",
	x"02", x"00", x"01", x"02", x"01", x"01", x"00", x"FF", x"FF", x"03", x"02", x"01",
	x"02", x"00", x"FF", x"01", x"01", x"FE", x"FF", x"FF", x"FC", x"FA", x"FC", x"FB",
	x"FE", x"00", x"FD", x"FD", x"00", x"02", x"00", x"03", x"04", x"01", x"02", x"FF",
	x"FD", x"FE", x"00", x"01", x"FF", x"00", x"FF", x"00", x"00", x"02", x"02", x"03",
	x"04", x"02", x"FE", x"FE", x"FE", x"FC", x"FC", x"FC", x"FA", x"FB", x"FE", x"FD",
	x"FE", x"01", x"00", x"01", x"02", x"02", x"FF", x"01", x"03", x"00", x"00", x"00",
	x"FF", x"01", x"03", x"02", x"00", x"02", x"01", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FA", x"F9", x"FB", x"FD", x"FF", x"FE", x"FE", x"00", x"00", x"01", x"02",
	x"03", x"05", x"03", x"02", x"00", x"FD", x"FE", x"FF", x"01", x"FE", x"FF", x"01",
	x"01", x"02", x"01", x"01", x"00", x"00", x"FD", x"FB", x"FC", x"FC", x"FD", x"FE",
	x"FD", x"FD", x"FF", x"02", x"02", x"01", x"01", x"01", x"02", x"01", x"FF", x"00",
	x"00", x"00", x"FD", x"FD", x"FD", x"FE", x"02", x"01", x"02", x"01", x"02", x"01",
	x"FF", x"00", x"00", x"00", x"FF", x"FD", x"FC", x"FC", x"FF", x"FE", x"FE", x"01",
	x"00", x"00", x"00", x"00", x"FF", x"01", x"02", x"FF", x"FE", x"FD", x"FD", x"FF",
	x"00", x"00", x"01", x"04", x"04", x"00", x"01", x"00", x"FF", x"FF", x"FD", x"FC",
	x"FB", x"FE", x"FF", x"FE", x"00", x"01", x"03", x"03", x"01", x"01", x"01", x"03",
	x"00", x"FB", x"FB", x"FD", x"FD", x"FF", x"FD", x"FD", x"FF", x"00", x"01", x"02",
	x"03", x"04", x"04", x"01", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE", x"FC", x"FD",
	x"FF", x"FF", x"01", x"02", x"03", x"03", x"01", x"FE", x"FD", x"FE", x"FE", x"FD",
	x"FC", x"FC", x"FD", x"00", x"00", x"00", x"01", x"01", x"03", x"01", x"00", x"01",
	x"01", x"00", x"FF", x"FE", x"FC", x"FE", x"01", x"01", x"00", x"01", x"00", x"01",
	x"02", x"FF", x"00", x"01", x"FD", x"FC", x"FB", x"FB", x"FC", x"FF", x"00", x"FF",
	x"FF", x"01", x"00", x"02", x"02", x"01", x"04", x"03", x"01", x"FD", x"FD", x"FF",
	x"FE", x"FF", x"FF", x"00", x"01", x"01", x"02", x"02", x"02", x"04", x"00", x"FE",
	x"FD", x"FB", x"FC", x"FD", x"FB", x"FA", x"FE", x"FF", x"FE", x"00", x"02", x"02",
	x"01", x"01", x"00", x"00", x"04", x"01", x"01", x"00", x"FE", x"00", x"01", x"03",
	x"00", x"01", x"03", x"FF", x"FE", x"FF", x"00", x"00", x"FE", x"FD", x"FB", x"F9",
	x"FC", x"FC", x"FD", x"FE", x"FE", x"00", x"01", x"00", x"FF", x"03", x"05", x"02",
	x"FF", x"01", x"02", x"01", x"03", x"01", x"00", x"04", x"03", x"02", x"00", x"00",
	x"00", x"FE", x"FE", x"F9", x"F9", x"FB", x"FB", x"FB", x"FA", x"FC", x"FF", x"00",
	x"02", x"02", x"02", x"04", x"03", x"02", x"01", x"00", x"01", x"01", x"02", x"00",
	x"FF", x"01", x"02", x"01", x"00", x"02", x"00", x"01", x"FF", x"FC", x"FC", x"FC",
	x"FF", x"FC", x"FC", x"FB", x"FB", x"FE", x"FE", x"FF", x"01", x"02", x"03", x"01",
	x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"02", x"02", x"03", x"04",
	x"03", x"04", x"02", x"01", x"FF", x"FF", x"FE", x"FA", x"F9", x"F9", x"FB", x"FB",
	x"FE", x"FD", x"FD", x"FF", x"FE", x"01", x"01", x"03", x"03", x"01", x"01", x"FF",
	x"FF", x"02", x"03", x"02", x"02", x"03", x"02", x"01", x"03", x"02", x"03", x"02",
	x"FC", x"FC", x"FB", x"FB", x"FA", x"FA", x"FA", x"FA", x"FD", x"FE", x"FF", x"00",
	x"03", x"04", x"02", x"02", x"01", x"02", x"01", x"00", x"FF", x"FE", x"00", x"01",
	x"01", x"03", x"02", x"02", x"03", x"02", x"FF", x"FD", x"00", x"00", x"FC", x"FB",
	x"FA", x"FB", x"FE", x"FD", x"FD", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"02",
	x"04", x"02", x"FF", x"FF", x"FF", x"01", x"00", x"FE", x"03", x"03", x"02", x"02",
	x"00", x"02", x"02", x"02", x"00", x"FD", x"FC", x"FB", x"FB", x"FB", x"FA", x"FC",
	x"FD", x"FE", x"FE", x"00", x"01", x"02", x"02", x"01", x"01", x"00", x"01", x"03",
	x"02", x"00", x"00", x"01", x"01", x"01", x"02", x"00", x"00", x"00", x"FC", x"FD",
	x"FD", x"FE", x"FE", x"FD", x"FD", x"FC", x"FE", x"FF", x"00", x"02", x"02", x"02",
	x"02", x"01", x"00", x"01", x"00", x"00", x"FF", x"FE", x"FF", x"FE", x"FD", x"FF",
	x"00", x"00", x"01", x"02", x"02", x"01", x"02", x"00", x"FF", x"00", x"FD", x"FD",
	x"FC", x"FE", x"FD", x"FE", x"01", x"FF", x"01", x"01", x"01", x"01", x"00", x"FE",
	x"FD", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"00", x"01", x"01", x"03",
	x"04", x"01", x"00", x"FE", x"FF", x"FD", x"FD", x"FE", x"FE", x"FF", x"FE", x"FE",
	x"FE", x"00", x"02", x"02", x"03", x"00", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE",
	x"FF", x"FE", x"FE", x"FF", x"01", x"03", x"03", x"03", x"00", x"FF", x"00", x"FF",
	x"FD", x"FB", x"FB", x"FD", x"00", x"FF", x"FF", x"04", x"03", x"04", x"01", x"01",
	x"02", x"01", x"01", x"FD", x"FC", x"FB", x"FA", x"FC", x"FC", x"FD", x"FE", x"00",
	x"02", x"FF", x"02", x"05", x"03", x"03", x"01", x"00", x"FE", x"FE", x"FF", x"FD",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"03", x"01", x"FF", x"00", x"FF",
	x"FD", x"FC", x"FD", x"FC", x"FD", x"00", x"FF", x"01", x"02", x"02", x"02", x"01",
	x"01", x"FF", x"FF", x"FF", x"FD", x"FD", x"FF", x"00", x"FE", x"FF", x"04", x"03",
	x"03", x"03", x"01", x"00", x"00", x"FE", x"FD", x"FE", x"FD", x"FB", x"FC", x"FC",
	x"FD", x"FF", x"01", x"01", x"FF", x"01", x"FF", x"00", x"01", x"00", x"01", x"00",
	x"00", x"FF", x"FE", x"00", x"00", x"02", x"02", x"02", x"03", x"01", x"03", x"02",
	x"FE", x"FF", x"FD", x"FB", x"FC", x"FA", x"FB", x"FC", x"FD", x"FE", x"FE", x"01",
	x"01", x"02", x"02", x"01", x"00", x"01", x"01", x"00", x"02", x"00", x"02", x"02",
	x"00", x"01", x"02", x"02", x"01", x"01", x"00", x"FD", x"FD", x"FC", x"FB", x"FD",
	x"FC", x"FC", x"FF", x"FE", x"FD", x"FE", x"00", x"02", x"02", x"02", x"00", x"01",
	x"01", x"00", x"FF", x"00", x"00", x"01", x"01", x"FF", x"01", x"01", x"04", x"03",
	x"FF", x"01", x"01", x"FF", x"FC", x"FB", x"FC", x"FB", x"FB", x"FB", x"FC", x"FF",
	x"01", x"FF", x"01", x"01", x"01", x"02", x"03", x"02", x"FF", x"01", x"FF", x"FE",
	x"FF", x"00", x"01", x"02", x"01", x"00", x"01", x"01", x"01", x"01", x"01", x"FF",
	x"FD", x"FE", x"FC", x"FB", x"FC", x"FE", x"FD", x"FC", x"FE", x"FF", x"01", x"01",
	x"02", x"01", x"01", x"02", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"04", x"04", x"02", x"01", x"01", x"00", x"00", x"FE", x"FD", x"FC", x"FC", x"FA",
	x"F9", x"FD", x"FD", x"FF", x"01", x"00", x"01", x"01", x"02", x"02", x"01", x"01",
	x"01", x"00", x"00", x"00", x"FF", x"00", x"01", x"02", x"02", x"01", x"01", x"00",
	x"00", x"FE", x"FE", x"FF", x"FE", x"FD", x"FC", x"FA", x"FB", x"FD", x"FD", x"FF",
	x"00", x"02", x"02", x"01", x"03", x"01", x"02", x"03", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"00", x"00", x"00", x"02", x"03", x"03", x"01", x"01", x"00", x"FE", x"FE",
	x"FD", x"FC", x"FC", x"FD", x"FD", x"FB", x"FE", x"FF", x"00", x"04", x"01", x"00",
	x"01", x"01", x"01", x"FF", x"01", x"02", x"01", x"02", x"FE", x"FF", x"01", x"01",
	x"01", x"00", x"01", x"00", x"00", x"FF", x"FD", x"FC", x"FD", x"FD", x"FC", x"FC",
	x"FD", x"FF", x"FF", x"00", x"02", x"01", x"04", x"03", x"01", x"02", x"01", x"FF",
	x"01", x"00", x"FE", x"FF", x"01", x"00", x"FE", x"01", x"00", x"00", x"01", x"FF",
	x"FE", x"FE", x"FE", x"FC", x"FD", x"FE", x"FE", x"00", x"01", x"00", x"00", x"01",
	x"02", x"02", x"01", x"01", x"02", x"00", x"FD", x"FD", x"FE", x"FF", x"FE", x"FD",
	x"FF", x"00", x"00", x"01", x"01", x"03", x"02", x"03", x"02", x"FE", x"FF", x"FE",
	x"FE", x"FD", x"FB", x"FC", x"FD", x"FF", x"FF", x"FF", x"01", x"01", x"02", x"01",
	x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"02", x"03", x"02", x"00", x"00",
	x"02", x"00", x"00", x"FF", x"FD", x"FF", x"FE", x"FC", x"FC", x"FC", x"FE", x"00",
	x"00", x"FF", x"00", x"04", x"02", x"02", x"01", x"01", x"01", x"00", x"FF", x"FD",
	x"FD", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"02", x"02", x"00", x"00", x"01",
	x"01", x"FF", x"FE", x"FD", x"FC", x"FD", x"FE", x"FE", x"00", x"02", x"02", x"02",
	x"02", x"01", x"01", x"02", x"FF", x"FC", x"FC", x"FD", x"FC", x"FD", x"FE", x"FD",
	x"00", x"02", x"02", x"02", x"03", x"04", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FE", x"FC", x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"02", x"02",
	x"01", x"00", x"FF", x"FF", x"FE", x"FD", x"FC", x"FE", x"00", x"FF", x"FE", x"00",
	x"02", x"02", x"03", x"02", x"01", x"02", x"01", x"FE", x"FD", x"FC", x"FD", x"FE",
	x"FC", x"FC", x"FD", x"00", x"00", x"FF", x"01", x"02", x"03", x"03", x"02", x"00",
	x"00", x"01", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FE", x"FF", x"01",
	x"01", x"FF", x"FD", x"FE", x"FC", x"FC", x"FD", x"FB", x"FD", x"FF", x"00", x"01",
	x"FF", x"02", x"04", x"04", x"02", x"00", x"03", x"01", x"FF", x"FF", x"FE", x"FF",
	x"00", x"00", x"FF", x"00", x"01", x"FF", x"00", x"FE", x"FD", x"FE", x"FE", x"FD",
	x"FC", x"FD", x"FC", x"FE", x"00", x"FF", x"02", x"01", x"02", x"02", x"01", x"01",
	x"01", x"01", x"01", x"00", x"FE", x"FD", x"FF", x"FF", x"FF", x"00", x"01", x"01",
	x"02", x"01", x"00", x"00", x"01", x"FE", x"FD", x"FD", x"FB", x"FB", x"FB", x"FC",
	x"FD", x"00", x"01", x"01", x"03", x"02", x"03", x"03", x"01", x"02", x"01", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"FE",
	x"FE", x"FC", x"FD", x"FC", x"FC", x"FD", x"FC", x"FF", x"FE", x"FE", x"01", x"03",
	x"03", x"02", x"01", x"00", x"01", x"02", x"02", x"00", x"FF", x"00", x"00", x"FD",
	x"FD", x"00", x"02", x"02", x"00", x"FF", x"01", x"01", x"FF", x"FD", x"FC", x"FB",
	x"FC", x"FC", x"FD", x"FD", x"FE", x"01", x"00", x"00", x"01", x"02", x"03", x"03",
	x"01", x"FF", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"01", x"00", x"00",
	x"01", x"02", x"00", x"FD", x"FC", x"FD", x"FD", x"FD", x"FC", x"FD", x"FE", x"FE",
	x"FE", x"FE", x"00", x"01", x"02", x"03", x"02", x"01", x"02", x"02", x"00", x"FF",
	x"00", x"01", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"01", x"FF", x"FE",
	x"FD", x"FD", x"FD", x"FC", x"FD", x"FE", x"FD", x"FE", x"FF", x"00", x"00", x"01",
	x"02", x"01", x"03", x"01", x"01", x"01", x"00", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"FF", x"FF", x"FE", x"FF", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FD",
	x"FE", x"FE", x"00", x"FF", x"FE", x"00", x"FF", x"01", x"03", x"01", x"01", x"00",
	x"00", x"FE", x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"02", x"02", x"02",
	x"02", x"00", x"FF", x"FF", x"FF", x"FE", x"FC", x"FD", x"FE", x"FD", x"FE", x"FF",
	x"00", x"01", x"02", x"01", x"FD", x"01", x"01", x"FF", x"00", x"FE", x"FE", x"FE",
	x"FF", x"FE", x"FF", x"03", x"02", x"03", x"02", x"01", x"01", x"02", x"01", x"FF",
	x"FF", x"FF", x"FD", x"FC", x"FB", x"FC", x"FE", x"FE", x"00", x"FF", x"00", x"01",
	x"01", x"03", x"00", x"02", x"FF", x"FF", x"FF", x"FC", x"FF", x"00", x"00", x"00",
	x"01", x"01", x"02", x"03", x"01", x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FE",
	x"FF", x"FF", x"FD", x"00", x"02", x"03", x"03", x"01", x"01", x"FF", x"FD", x"FD",
	x"FD", x"FF", x"FD", x"FD", x"FD", x"FC", x"FF", x"01", x"03", x"03", x"02", x"03",
	x"04", x"03", x"01", x"00", x"00", x"FE", x"FD", x"FC", x"FD", x"FE", x"FF", x"00",
	x"00", x"00", x"00", x"01", x"01", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FF",
	x"FF", x"01", x"01", x"00", x"01", x"02", x"03", x"03", x"02", x"01", x"00", x"00",
	x"FE", x"FC", x"FE", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"01",
	x"01", x"02", x"02", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"00",
	x"FF", x"00", x"02", x"03", x"02", x"00", x"FF", x"FE", x"FD", x"FD", x"FB", x"FB",
	x"FC", x"FB", x"FB", x"FD", x"00", x"02", x"03", x"02", x"02", x"03", x"02", x"03",
	x"03", x"03", x"02", x"FF", x"FF", x"FE", x"FE", x"00", x"00", x"FF", x"FE", x"FD",
	x"FD", x"FD", x"FE", x"FE", x"FF", x"FE", x"FE", x"FD", x"FD", x"FD", x"FF", x"01",
	x"00", x"01", x"02", x"04", x"04", x"02", x"02", x"01", x"01", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FE", x"FE", x"00", x"02", x"02", x"00", x"FF", x"00", x"FF",
	x"FE", x"FC", x"FD", x"FD", x"FE", x"FD", x"FC", x"FE", x"00", x"01", x"03", x"04",
	x"02", x"02", x"02", x"FF", x"FF", x"00", x"00", x"01", x"00", x"FD", x"FD", x"00",
	x"01", x"00", x"01", x"01", x"00", x"00", x"FE", x"FD", x"FD", x"FE", x"FE", x"FB",
	x"FA", x"FB", x"FE", x"00", x"00", x"01", x"02", x"04", x"04", x"04", x"03", x"03",
	x"00", x"FE", x"FF", x"FD", x"FE", x"01", x"FF", x"FD", x"FE", x"FF", x"FF", x"01",
	x"02", x"FF", x"00", x"FE", x"FC", x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"FD",
	x"00", x"02", x"03", x"03", x"01", x"02", x"00", x"00", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"FD", x"FF", x"00", x"FF", x"02", x"00", x"00", x"01", x"01", x"FF", x"FE",
	x"FE", x"FD", x"FC", x"FD", x"FC", x"FD", x"00", x"00", x"00", x"01", x"02", x"01",
	x"02", x"02", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FE", x"FD", x"FD", x"FC", x"FC", x"FE",
	x"01", x"02", x"01", x"01", x"02", x"01", x"02", x"01", x"01", x"02", x"02", x"00",
	x"FC", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"00", x"FF", x"FF", x"01",
	x"00", x"00", x"FE", x"FE", x"FE", x"FF", x"00", x"FE", x"FE", x"00", x"02", x"03",
	x"02", x"01", x"01", x"00", x"00", x"FE", x"FE", x"FF", x"FF", x"FF", x"FD", x"FD",
	x"FE", x"00", x"02", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"FF",
	x"00", x"00", x"FF", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"00",
	x"02", x"03", x"01", x"01", x"01", x"00", x"FF", x"FD", x"FD", x"FD", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"01", x"02", x"02", x"02", x"02", x"00", x"FE", x"FE", x"FD",
	x"FF", x"00", x"FE", x"FD", x"FD", x"FF", x"00", x"00", x"02", x"02", x"02", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"FE", x"FD", x"FE", x"FF", x"FF", x"01", x"00",
	x"00", x"01", x"00", x"01", x"01", x"00", x"FF", x"FE", x"FD", x"FC", x"FE", x"FF",
	x"FF", x"01", x"FF", x"00", x"02", x"01", x"01", x"01", x"01", x"FF", x"FD", x"FE",
	x"FD", x"FF", x"01", x"FF", x"00", x"00", x"00", x"01", x"02", x"01", x"01", x"01",
	x"FF", x"FC", x"FD", x"FC", x"FD", x"FD", x"FD", x"FE", x"FF", x"01", x"01", x"01",
	x"02", x"04", x"04", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FD", x"FC", x"FF",
	x"FE", x"FF", x"00", x"FF", x"01", x"02", x"00", x"FF", x"FF", x"FF", x"FE", x"FD",
	x"FD", x"FC", x"00", x"01", x"01", x"01", x"02", x"03", x"01", x"01", x"FF", x"00",
	x"01", x"00", x"FF", x"FC", x"FE", x"FF", x"FF", x"01", x"01", x"01", x"00", x"01",
	x"FF", x"FD", x"FF", x"FE", x"FE", x"FD", x"FC", x"FC", x"FE", x"FF", x"00", x"01",
	x"02", x"01", x"01", x"03", x"03", x"01", x"02", x"02", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FD", x"00", x"01", x"00", x"01", x"00", x"FF", x"FC", x"FD",
	x"FD", x"FC", x"FE", x"FE", x"FE", x"FF", x"01", x"02", x"03", x"05", x"05", x"04",
	x"03", x"01", x"00", x"01", x"FF", x"FE", x"FE", x"FE", x"FC", x"FC", x"FD", x"FD",
	x"FE", x"00", x"00", x"FF", x"FE", x"FF", x"FD", x"FF", x"FF", x"FE", x"00", x"00",
	x"00", x"00", x"01", x"03", x"02", x"03", x"03", x"01", x"01", x"01", x"01", x"FE",
	x"FD", x"FD", x"FC", x"FE", x"FE", x"FE", x"00", x"01", x"00", x"FF", x"00", x"01",
	x"01", x"00", x"FD", x"FB", x"FB", x"FD", x"FE", x"FE", x"00", x"00", x"00", x"01",
	x"02", x"02", x"04", x"05", x"03", x"01", x"00", x"FF", x"FF", x"00", x"FF", x"FD",
	x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"FD", x"FD", x"FE", x"FF",
	x"FF", x"FE", x"FD", x"FF", x"01", x"02", x"02", x"02", x"04", x"05", x"04", x"02",
	x"03", x"02", x"00", x"FF", x"FC", x"FB", x"FD", x"FD", x"FD", x"FE", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FF", x"FE", x"FE", x"FF", x"00",
	x"01", x"01", x"02", x"02", x"02", x"02", x"01", x"02", x"01", x"00", x"00", x"FE",
	x"FE", x"FE", x"FE", x"00", x"00", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"FE", x"FF", x"FE", x"FD", x"FC", x"FD", x"FE", x"00", x"00", x"00", x"03", x"04",
	x"05", x"04", x"03", x"02", x"02", x"01", x"00", x"FE", x"FE", x"FE", x"FE", x"FC",
	x"FB", x"FF", x"00", x"FF", x"FF", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FF",
	x"FE", x"00", x"00", x"00", x"02", x"05", x"05", x"03", x"02", x"00", x"01", x"02",
	x"FF", x"FF", x"FD", x"FD", x"FD", x"FC", x"FD", x"FC", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"02", x"01", x"00", x"00", x"FD", x"00", x"FF", x"FF", x"00", x"FF", x"01",
	x"00", x"01", x"01", x"00", x"02", x"02", x"01", x"FF", x"FF", x"FE", x"FE", x"00",
	x"FE", x"FE", x"00", x"00", x"00", x"FF", x"00", x"01", x"02", x"01", x"FD", x"FC",
	x"FD", x"FD", x"FD", x"FD", x"FF", x"FE", x"FF", x"00", x"FF", x"02", x"04", x"03",
	x"02", x"01", x"01", x"00", x"00", x"FF", x"FD", x"FF", x"FD", x"FC", x"FE", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"02", x"02", x"FF", x"FE", x"FE", x"FD", x"FC",
	x"FE", x"FF", x"00", x"01", x"00", x"00", x"00", x"03", x"02", x"02", x"01", x"FE",
	x"FE", x"FE", x"FE", x"FC", x"FE", x"01", x"FF", x"FF", x"FF", x"FF", x"02", x"02",
	x"01", x"FF", x"01", x"01", x"FF", x"FF", x"FD", x"FD", x"FF", x"FF", x"FF", x"FE",
	x"01", x"01", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FD", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"01", x"01", x"03", x"01", x"00", x"01", x"01", x"00", x"FE",
	x"FE", x"FD", x"FD", x"FE", x"FD", x"FD", x"00", x"01", x"03", x"03", x"00", x"00",
	x"01", x"00", x"FE", x"FD", x"FE", x"FE", x"FD", x"FD", x"FD", x"FF", x"01", x"02",
	x"02", x"01", x"02", x"02", x"02", x"02", x"01", x"01", x"00", x"00", x"FE", x"FD",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FE", x"00", x"01", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"02", x"03", x"04", x"03", x"02",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FD", x"FE", x"FF", x"00",
	x"01", x"FF", x"FE", x"FE", x"FF", x"FC", x"FB", x"FE", x"FD", x"FE", x"FF", x"FE",
	x"00", x"02", x"04", x"03", x"03", x"05", x"04", x"03", x"01", x"FF", x"FF", x"FE",
	x"FE", x"FD", x"FC", x"FD", x"FD", x"FF", x"FF", x"FD", x"FF", x"01", x"01", x"FE",
	x"FE", x"FF", x"FD", x"FE", x"FD", x"FD", x"FE", x"02", x"03", x"01", x"02", x"03",
	x"04", x"05", x"03", x"01", x"00", x"00", x"FD", x"FB", x"FD", x"FE", x"FF", x"FF",
	x"FE", x"FD", x"FE", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FE", x"FD", x"FD",
	x"FE", x"00", x"FE", x"00", x"01", x"02", x"03", x"04", x"03", x"01", x"03", x"03",
	x"01", x"00", x"FD", x"FD", x"FE", x"FE", x"FD", x"FD", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FD", x"FB", x"FC", x"FB", x"FC", x"FE", x"FE", x"02",
	x"03", x"03", x"03", x"04", x"05", x"03", x"03", x"02", x"01", x"00", x"FF", x"FE",
	x"FB", x"FC", x"FD", x"FD", x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE",
	x"FE", x"FF", x"FE", x"FE", x"FF", x"00", x"02", x"02", x"01", x"03", x"03", x"03",
	x"02", x"01", x"02", x"01", x"00", x"FE", x"FD", x"FE", x"FD", x"FD", x"FD", x"FE",
	x"FF", x"00", x"02", x"00", x"00", x"00", x"FE", x"FD", x"FD", x"FD", x"FE", x"00",
	x"FE", x"FE", x"00", x"01", x"02", x"03", x"03", x"03", x"02", x"02", x"00", x"FF",
	x"01", x"00", x"00", x"FE", x"FD", x"FF", x"FF", x"00", x"FF", x"FE", x"FE", x"FF",
	x"FE", x"FC", x"FD", x"FD", x"FE", x"FF", x"FD", x"FD", x"01", x"02", x"01", x"02",
	x"03", x"04", x"05", x"04", x"02", x"00", x"01", x"FF", x"FD", x"FD", x"FD", x"FD",
	x"FE", x"FD", x"FD", x"FE", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FE", x"FE", x"00", x"01", x"01", x"01", x"02", x"01", x"02", x"03", x"00", x"01",
	x"01", x"FF", x"FD", x"FD", x"FD", x"FD", x"FF", x"FF", x"FD", x"FF", x"00", x"00",
	x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"00", x"FF", x"FD", x"FD", x"FD",
	x"FE", x"FF", x"00", x"01", x"01", x"01", x"03", x"01", x"01", x"02", x"FF", x"FF",
	x"FF", x"FD", x"FE", x"FF", x"00", x"00", x"00", x"01", x"FF", x"00", x"00", x"FF",
	x"FE", x"FF", x"FF", x"FC", x"FD", x"FE", x"FE", x"FF", x"01", x"01", x"02", x"03",
	x"04", x"02", x"01", x"01", x"01", x"01", x"00", x"FE", x"FB", x"FD", x"FC", x"FB",
	x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"03", x"02", x"01", x"01", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"01", x"01", x"01", x"00",
	x"00", x"FD", x"FE", x"00", x"FE", x"FD", x"FD", x"FE", x"FF", x"00", x"01", x"01",
	x"03", x"02", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FD", x"FF", x"FF",
	x"00", x"00", x"01", x"02", x"00", x"00", x"FF", x"00", x"01", x"FF", x"FE", x"FD",
	x"FE", x"FE", x"FD", x"FF", x"FF", x"FF", x"01", x"01", x"01", x"01", x"03", x"01",
	x"FF", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"02", x"02",
	x"01", x"02", x"00", x"FF", x"FC", x"FC", x"FE", x"FC", x"FD", x"FD", x"FD", x"FF",
	x"00", x"01", x"01", x"03", x"04", x"02", x"02", x"01", x"00", x"FF", x"00", x"FF",
	x"FE", x"00", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"FE", x"FF", x"FE",
	x"FD", x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"03", x"03", x"02", x"03",
	x"02", x"01", x"00", x"FF", x"FE", x"FD", x"FC", x"FC", x"FD", x"FE", x"FF", x"01",
	x"00", x"01", x"01", x"00", x"01", x"01", x"FF", x"FE", x"FE", x"FC", x"FC", x"FE",
	x"FF", x"00", x"02", x"01", x"02", x"02", x"01", x"01", x"03", x"02", x"00", x"FF",
	x"FF", x"FD", x"FD", x"FE", x"FD", x"FD", x"FF", x"00", x"FF", x"FF", x"00", x"00",
	x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FF", x"FF", x"01", x"02",
	x"01", x"03", x"03", x"03", x"00", x"00", x"01", x"FF", x"FF", x"FD", x"FC", x"FE",
	x"FE", x"FD", x"FE", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FE",
	x"FE", x"FF", x"FE", x"FE", x"FF", x"00", x"02", x"03", x"03", x"02", x"02", x"02",
	x"01", x"01", x"00", x"FF", x"FE", x"FD", x"FE", x"FC", x"FD", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"00", x"01", x"00", x"FE", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"01", x"01", x"01", x"04", x"05", x"04", x"02", x"00", x"00", x"FE", x"FF",
	x"FE", x"FD", x"FE", x"FC", x"FC", x"FC", x"FE", x"00", x"00", x"01", x"FE", x"FE",
	x"FF", x"FE", x"FF", x"FE", x"00", x"FF", x"FF", x"01", x"00", x"02", x"02", x"03",
	x"02", x"01", x"02", x"01", x"01", x"00", x"FE", x"FD", x"FD", x"FE", x"FC", x"FD",
	x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"01", x"01", x"FE", x"FE", x"FD", x"FD",
	x"FF", x"FE", x"00", x"01", x"03", x"03", x"02", x"03", x"02", x"02", x"02", x"02",
	x"00", x"FE", x"FE", x"FD", x"FC", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"00", x"FF", x"FF", x"FF", x"FD", x"FD", x"FE", x"00", x"FF", x"00", x"04", x"01",
	x"02", x"03", x"03", x"04", x"03", x"02", x"FF", x"00", x"00", x"FD", x"FE", x"FC",
	x"FB", x"FB", x"FC", x"FE", x"FE", x"01", x"02", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FE", x"FE", x"FD", x"FE", x"FF", x"02", x"02", x"01", x"03", x"01",
	x"00", x"02", x"00", x"FF", x"FF", x"FF", x"FD", x"FE", x"FF", x"FD", x"00", x"01",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FD", x"FE", x"FF", x"FE", x"FD",
	x"FE", x"00", x"00", x"00", x"00", x"01", x"03", x"04", x"03", x"01", x"02", x"01",
	x"FF", x"FF", x"FD", x"FE", x"FF", x"FE", x"FD", x"FC", x"FF", x"00", x"00", x"01",
	x"FE", x"FE", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"01",
	x"03", x"04", x"03", x"02", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FC", x"FD", x"FE", x"FF", x"00", x"FF", x"FF", x"01", x"02", x"01", x"01", x"01",
	x"FF", x"FE", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"01",
	x"02", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"01", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF",
	x"FF", x"00", x"01", x"01", x"01", x"03", x"02", x"01", x"02", x"01", x"FF", x"FE",
	x"FE", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"02", x"02",
	x"01", x"01", x"FF", x"FF", x"FE", x"FE", x"FD", x"FC", x"FE", x"00", x"00", x"01",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FE", x"FE", x"FD", x"FC", x"FF",
	x"01", x"04", x"02", x"01", x"02", x"02", x"02", x"01", x"01", x"FF", x"FE", x"FE",
	x"FB", x"FA", x"FD", x"FF", x"FF", x"FD", x"FE", x"FF", x"01", x"01", x"FE", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"01", x"00", x"01", x"03", x"04",
	x"03", x"01", x"FF", x"FF", x"FF", x"FD", x"FC", x"FB", x"FB", x"FC", x"FB", x"FC",
	x"FD", x"00", x"04", x"03", x"02", x"02", x"02", x"01", x"00", x"00", x"FE", x"FE",
	x"FF", x"FD", x"FD", x"FF", x"00", x"01", x"03", x"04", x"01", x"02", x"02", x"FF",
	x"FF", x"00", x"FF", x"FD", x"FE", x"FD", x"FC", x"FE", x"FE", x"FF", x"00", x"00",
	x"FF", x"FE", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"00",
	x"03", x"02", x"01", x"03", x"03", x"03", x"01", x"01", x"FE", x"FC", x"FD", x"FC",
	x"FD", x"FE", x"FD", x"FC", x"FE", x"FF", x"FF", x"01", x"01", x"00", x"00", x"FF",
	x"FE", x"FD", x"00", x"00", x"00", x"00", x"FF", x"00", x"03", x"03", x"03", x"01",
	x"02", x"02", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FC", x"FB", x"FE", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"00", x"01", x"FF", x"FF", x"00", x"00", x"FF", x"FE",
	x"FE", x"FF", x"02", x"03", x"01", x"01", x"03", x"04", x"03", x"01", x"00", x"00",
	x"FF", x"FE", x"FC", x"FB", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FE", x"FF", x"00", x"FF", x"FE", x"FE", x"FE", x"00", x"01", x"02", x"02", x"02",
	x"03", x"03", x"03", x"02", x"01", x"00", x"FF", x"FE", x"FD", x"FD", x"FE", x"FE",
	x"FE", x"FD", x"FD", x"FE", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF",
	x"00", x"00", x"FF", x"FD", x"FE", x"01", x"02", x"02", x"03", x"03", x"02", x"01",
	x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FC", x"FD", x"FE", x"FF", x"01", x"00",
	x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE", x"FD", x"FF", x"00",
	x"00", x"01", x"01", x"02", x"02", x"03", x"02", x"00", x"01", x"00", x"FF", x"FE",
	x"FE", x"FE", x"FD", x"FF", x"FD", x"FE", x"FF", x"01", x"02", x"01", x"02", x"02",
	x"00", x"FF", x"FD", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"01",
	x"01", x"02", x"03", x"02", x"00", x"FF", x"FF", x"FF", x"01", x"00", x"FE", x"FE",
	x"FF", x"00", x"00", x"01", x"00", x"00", x"01", x"FF", x"FD", x"FD", x"FE", x"FF",
	x"FD", x"FD", x"FE", x"00", x"01", x"01", x"01", x"00", x"01", x"02", x"01", x"02",
	x"01", x"01", x"00", x"FE", x"FC", x"FD", x"FF", x"FE", x"FF", x"FF", x"FE", x"00",
	x"01", x"02", x"02", x"02", x"00", x"FE", x"FE", x"FD", x"FC", x"FF", x"00", x"FF",
	x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"00", x"FF", x"01", x"01", x"01", x"00", x"00", x"02", x"00", x"FF",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FC", x"FE", x"FF", x"FD", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"01", x"02", x"FF", x"FF", x"00", x"00", x"FF", x"01",
	x"02", x"02", x"02", x"01", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FC", x"FB",
	x"FD", x"FE", x"FF", x"00", x"02", x"01", x"01", x"02", x"00", x"00", x"02", x"00",
	x"FE", x"FD", x"FD", x"FE", x"FE", x"00", x"FF", x"00", x"02", x"02", x"01", x"02",
	x"03", x"01", x"00", x"00", x"FF", x"FF", x"00", x"FE", x"FC", x"FB", x"FC", x"FC",
	x"FE", x"FF", x"FF", x"01", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"01", x"00",
	x"FF", x"01", x"03", x"03", x"03", x"04", x"03", x"02", x"01", x"FF", x"FD", x"FD",
	x"FD", x"FC", x"FB", x"FB", x"FC", x"FC", x"FE", x"FF", x"FF", x"01", x"03", x"01",
	x"01", x"02", x"00", x"00", x"01", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01",
	x"01", x"02", x"02", x"00", x"00", x"01", x"FF", x"FD", x"FC", x"FC", x"FC", x"FD",
	x"FE", x"FD", x"FE", x"FF", x"01", x"01", x"02", x"03", x"03", x"01", x"00", x"FE",
	x"FD", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"01", x"02", x"02", x"04", x"03",
	x"02", x"FF", x"00", x"FF", x"FE", x"FE", x"FC", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"00", x"FF", x"FE", x"FF", x"FF", x"01", x"01", x"01", x"00", x"FF", x"01", x"01",
	x"01", x"02", x"03", x"03", x"01", x"01", x"00", x"00", x"02", x"00", x"FE", x"FC",
	x"FB", x"FB", x"FC", x"FD", x"FC", x"FF", x"FF", x"00", x"01", x"00", x"02", x"02",
	x"02", x"01", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"02", x"01",
	x"00", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FD", x"FD", x"FC", x"FD", x"FE",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"01", x"FF", x"FF", x"FE", x"FF", x"00",
	x"00", x"00", x"FF", x"01", x"01", x"01", x"02", x"02", x"04", x"02", x"01", x"FF",
	x"FE", x"FF", x"FE", x"FD", x"FB", x"FB", x"FC", x"FC", x"FF", x"FF", x"00", x"02",
	x"01", x"00", x"FF", x"00", x"01", x"FF", x"00", x"FF", x"FF", x"01", x"01", x"02",
	x"02", x"02", x"01", x"02", x"02", x"00", x"00", x"FE", x"FD", x"FC", x"FB", x"FC",
	x"FD", x"FE", x"FD", x"FE", x"FF", x"00", x"01", x"01", x"03", x"03", x"01", x"01",
	x"00", x"FF", x"00", x"00", x"FE", x"FE", x"FF", x"00", x"FF", x"00", x"00", x"02",
	x"02", x"01", x"FF", x"FF", x"FF", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"00",
	x"FE", x"00", x"02", x"02", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FD", x"FF",
	x"00", x"FF", x"FF", x"00", x"01", x"01", x"02", x"01", x"FF", x"01", x"01", x"FF",
	x"FF", x"FD", x"FD", x"FE", x"FF", x"FD", x"FE", x"00", x"00", x"FF", x"FE", x"00",
	x"01", x"02", x"03", x"01", x"FF", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"00",
	x"00", x"FF", x"00", x"01", x"01", x"00", x"00", x"FF", x"FD", x"FF", x"FF", x"FD",
	x"FE", x"00", x"00", x"00", x"01", x"00", x"FF", x"01", x"00", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FD", x"FE", x"01", x"01", x"00", x"00", x"01", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"00", x"01", x"01", x"01", x"02", x"00", x"00", x"01", x"00", x"FE", x"FD", x"FE",
	x"FD", x"FD", x"FF", x"00", x"00", x"01", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FE", x"00", x"00", x"01", x"02", x"00", x"00", x"01", x"00",
	x"00", x"FE", x"FF", x"FE", x"FE", x"FE", x"FD", x"FF", x"00", x"FF", x"FE", x"FF",
	x"00", x"01", x"02", x"00", x"FE", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"FF", x"01", x"02", x"03", x"03", x"01", x"00", x"FF", x"FE", x"FE", x"FC",
	x"FB", x"FC", x"FE", x"FD", x"FC", x"FF", x"00", x"01", x"02", x"01", x"02", x"02",
	x"01", x"00", x"FF", x"FE", x"FF", x"00", x"FF", x"FF", x"FF", x"01", x"03", x"01",
	x"02", x"03", x"02", x"01", x"FF", x"FE", x"FD", x"FD", x"FE", x"FC", x"FB", x"FC",
	x"FD", x"FD", x"FD", x"FF", x"FF", x"01", x"02", x"01", x"03", x"02", x"01", x"01",
	x"00", x"01", x"01", x"02", x"02", x"02", x"01", x"00", x"01", x"00", x"00", x"FE",
	x"FD", x"FD", x"FB", x"FA", x"FB", x"FC", x"FD", x"FE", x"00", x"FF", x"00", x"03",
	x"02", x"02", x"02", x"02", x"01", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00",
	x"01", x"01", x"00", x"01", x"00", x"00", x"01", x"FF", x"FF", x"FF", x"FE", x"FD",
	x"FC", x"FC", x"FC", x"FD", x"FD", x"FE", x"FF", x"00", x"01", x"00", x"01", x"02",
	x"00", x"00", x"01", x"00", x"00", x"00", x"01", x"01", x"02", x"03", x"02", x"02",
	x"02", x"00", x"FF", x"FE", x"FE", x"FD", x"FD", x"FB", x"FA", x"FC", x"FC", x"FD",
	x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"02", x"02", x"01", x"01", x"01",
	x"02", x"03", x"03", x"02", x"01", x"02", x"01", x"00", x"00", x"FF", x"FD", x"FC",
	x"FC", x"FB", x"FB", x"FD", x"FD", x"FD", x"FC", x"FD", x"FF", x"02", x"02", x"01",
	x"02", x"02", x"01", x"00", x"01", x"00", x"00", x"00", x"FF", x"FE", x"00", x"02",
	x"02", x"02", x"02", x"02", x"01", x"00", x"FF", x"FE", x"FE", x"FD", x"FC", x"FC",
	x"FD", x"FD", x"FC", x"FE", x"FF", x"FF", x"00", x"01", x"00", x"00", x"01", x"00",
	x"FF", x"01", x"01", x"02", x"03", x"02", x"02", x"02", x"03", x"02", x"02", x"02",
	x"00", x"FF", x"FE", x"FC", x"FB", x"FA", x"FB", x"FA", x"FB", x"FC", x"FD", x"FF",
	x"01", x"01", x"01", x"03", x"04", x"02", x"01", x"00", x"FF", x"FF", x"00", x"01",
	x"00", x"02", x"02", x"00", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FC", x"FD",
	x"FC", x"FC", x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"02", x"01", x"01",
	x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"02",
	x"01", x"01", x"02", x"00", x"00", x"01", x"00", x"FF", x"FE", x"FC", x"FC", x"FD",
	x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"FE",
	x"FE", x"FE", x"FF", x"00", x"02", x"01", x"01", x"03", x"02", x"00", x"00", x"00",
	x"FF", x"FE", x"FE", x"FD", x"FD", x"FE", x"FD", x"FD", x"FF", x"00", x"00", x"00",
	x"01", x"00", x"01", x"02", x"00", x"FF", x"00", x"01", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"01", x"01", x"FF", x"FE", x"FF", x"FF", x"00", x"00",
	x"FE", x"FE", x"00", x"FF", x"FF", x"01", x"03", x"02", x"01", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FE", x"00", x"FF", x"00", x"02", x"01",
	x"00", x"00", x"02", x"01", x"00", x"FF", x"FE", x"FE", x"FF", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"00", x"02", x"02", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FD", x"FD", x"FE", x"FE", x"FE", x"00", x"00", x"01", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"02", x"02", x"01", x"01",
	x"01", x"01", x"00", x"FE", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FD",
	x"FF", x"FF", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"01", x"02", x"02", x"01", x"01", x"02", x"01", x"01", x"00",
	x"FE", x"FC", x"FB", x"FA", x"FA", x"FC", x"FD", x"FE", x"FF", x"FF", x"00", x"01",
	x"03", x"03", x"02", x"02", x"00", x"FF", x"00", x"00", x"FF", x"00", x"01", x"01",
	x"00", x"01", x"01", x"02", x"02", x"00", x"FE", x"FE", x"FE", x"FD", x"FC", x"FB",
	x"FD", x"FD", x"FE", x"FE", x"FE", x"00", x"01", x"00", x"00", x"00", x"02", x"02",
	x"02", x"01", x"00", x"01", x"00", x"00", x"01", x"01", x"01", x"03", x"02", x"00",
	x"FF", x"00", x"FF", x"FD", x"FD", x"FC", x"FB", x"FB", x"FC", x"FC", x"FE", x"00",
	x"01", x"02", x"01", x"01", x"01", x"02", x"02", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"01", x"02", x"02", x"02", x"01", x"01", x"02", x"01", x"00", x"FF", x"FD",
	x"FC", x"FC", x"FC", x"FB", x"FD", x"FD", x"FC", x"FC", x"FE", x"00", x"01", x"01",
	x"01", x"00", x"FF", x"01", x"02", x"01", x"03", x"02", x"01", x"01", x"01", x"02",
	x"03", x"03", x"01", x"FF", x"FE", x"FD", x"FC", x"FD", x"FC", x"FB", x"FB", x"FC",
	x"FC", x"FE", x"00", x"FF", x"01", x"01", x"00", x"01", x"02", x"02", x"FF", x"FF",
	x"00", x"00", x"01", x"02", x"02", x"01", x"02", x"02", x"00", x"01", x"01", x"FF",
	x"FE", x"FD", x"FD", x"FB", x"FC", x"FD", x"FC", x"FD", x"FE", x"FE", x"FF", x"01",
	x"00", x"01", x"03", x"02", x"01", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"03", x"02", x"01", x"01", x"01", x"02", x"02", x"00", x"FF", x"FD", x"FD", x"FB",
	x"FA", x"FC", x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"02", x"02", x"01", x"01",
	x"01", x"00", x"00", x"00", x"00", x"02", x"02", x"00", x"01", x"02", x"02", x"02",
	x"01", x"FF", x"FD", x"FE", x"FE", x"FD", x"FC", x"FB", x"FC", x"FC", x"FC", x"FD",
	x"FF", x"02", x"03", x"01", x"01", x"02", x"02", x"03", x"02", x"00", x"FF", x"FF",
	x"FE", x"FD", x"FE", x"00", x"01", x"00", x"00", x"FF", x"01", x"01", x"00", x"FF",
	x"FF", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"01",
	x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"01", x"00", x"02", x"03", x"02", x"00", x"00", x"FF", x"FE", x"FE", x"FD", x"FE",
	x"FD", x"FC", x"FC", x"FD", x"FF", x"01", x"01", x"02", x"01", x"00", x"00", x"00",
	x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"01", x"01", x"01", x"01", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FD", x"FD", x"FE", x"FE", x"FE", x"FF", x"00", x"01",
	x"01", x"00", x"00", x"01", x"02", x"02", x"00", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FD", x"FF", x"01", x"01", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"00", x"00", x"FF", x"00", x"00", x"01", x"02", x"02", x"01",
	x"00", x"00", x"FE", x"FE", x"FD", x"FC", x"FD", x"FF", x"00", x"FF", x"00", x"01",
	x"01", x"02", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FE", x"FF", x"FF",
	x"FE", x"FE", x"00", x"02", x"02", x"00", x"01", x"01", x"01", x"01", x"00", x"00",
	x"00", x"FF", x"FD", x"FC", x"FE", x"FF", x"00", x"00", x"FF", x"FE", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"02", x"02", x"02",
	x"01", x"02", x"02", x"02", x"00", x"FD", x"FD", x"FB", x"FB", x"FC", x"FD", x"FE",
	x"FD", x"FF", x"00", x"00", x"02", x"03", x"02", x"02", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FE", x"FE", x"00", x"01", x"01", x"00", x"01", x"00", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FD", x"FB", x"FC", x"FD", x"FD", x"FF", x"00", x"01",
	x"01", x"02", x"02", x"01", x"01", x"02", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"FF", x"FF", x"00", x"FE", x"FD",
	x"FD", x"FD", x"FE", x"FE", x"00", x"FF", x"FE", x"00", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"02", x"01", x"01", x"00", x"FF", x"01", x"02",
	x"03", x"01", x"00", x"FF", x"FD", x"FD", x"FC", x"FC", x"FC", x"FD", x"FD", x"FC",
	x"FC", x"00", x"02", x"02", x"02", x"02", x"01", x"02", x"01", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"01", x"02", x"01", x"00", x"00", x"00", x"FF", x"FF",
	x"FE", x"FD", x"FC", x"FC", x"FC", x"FD", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"00", x"01", x"02", x"02", x"01", x"01", x"00", x"01", x"00", x"00", x"01", x"02",
	x"02", x"01", x"01", x"00", x"FF", x"00", x"FF", x"FD", x"FC", x"FC", x"FA", x"FB",
	x"FC", x"FE", x"FE", x"FF", x"00", x"01", x"02", x"01", x"03", x"04", x"02", x"00",
	x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"01", x"02", x"02", x"02", x"01",
	x"01", x"FE", x"FC", x"FC", x"FD", x"FE", x"FC", x"FB", x"FC", x"FD", x"FE", x"FF",
	x"02", x"02", x"01", x"01", x"01", x"01", x"02", x"02", x"02", x"01", x"FF", x"FD",
	x"FE", x"00", x"01", x"02", x"01", x"01", x"00", x"01", x"00", x"FF", x"FF", x"FD",
	x"FD", x"FB", x"F9", x"FC", x"FD", x"FE", x"FF", x"FF", x"01", x"02", x"03", x"03",
	x"02", x"01", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"02", x"02", x"01", x"00", x"FE", x"FD", x"FE", x"FE", x"FD", x"FD", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"01", x"02", x"02", x"02", x"01", x"02", x"01", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"02", x"02", x"02", x"01",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE", x"FD", x"FE", x"FF", x"00",
	x"01", x"00", x"FF", x"00", x"01", x"00", x"FF", x"FE", x"FE", x"00", x"00", x"02",
	x"02", x"02", x"02", x"01", x"01", x"00", x"00", x"01", x"00", x"FE", x"FC", x"FC",
	x"FD", x"FE", x"FE", x"FD", x"FD", x"FF", x"FF", x"00", x"00", x"01", x"02", x"02",
	x"02", x"FF", x"FF", x"00", x"01", x"FF", x"FE", x"FF", x"00", x"01", x"00", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FE", x"FE", x"FF", x"01",
	x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FD", x"FF", x"01", x"01", x"00", x"01", x"02", x"01", x"00", x"00", x"01",
	x"01", x"01", x"FF", x"FE", x"FD", x"FD", x"FE", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"00", x"01", x"00", x"FF", x"FF", x"FE", x"FD", x"FE", x"FE", x"FF", x"01",
	x"00", x"00", x"01", x"03", x"03", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FF",
	x"FE", x"FF", x"FE", x"FE", x"00", x"01", x"02", x"02", x"01", x"00", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"FE", x"FD", x"FE", x"FE", x"FD", x"FF", x"00", x"00", x"01",
	x"01", x"00", x"01", x"02", x"01", x"00", x"00", x"00", x"FF", x"00", x"00", x"01",
	x"00", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FD", x"FC", x"FB", x"FB", x"FD",
	x"FD", x"FD", x"FF", x"00", x"01", x"03", x"04", x"03", x"03", x"04", x"03", x"01",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"FD", x"FE", x"00", x"FF", x"FE", x"FE", x"00",
	x"01", x"00", x"00", x"FE", x"FE", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"02", x"03", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"FF", x"FE", x"FF", x"FE",
	x"FD", x"FC", x"FC", x"FC", x"FD", x"FF", x"00", x"00", x"01", x"01", x"01", x"00",
	x"01", x"01", x"01", x"00", x"FF", x"00", x"00", x"01", x"01", x"02", x"02", x"01",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FD", x"FD", x"FC", x"FB", x"FC", x"FC",
	x"FD", x"FF", x"00", x"01", x"01", x"03", x"03", x"02", x"03", x"03", x"02", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"00", x"00", x"01",
	x"02", x"02", x"00", x"00", x"FF", x"00", x"01", x"00", x"01", x"01", x"00", x"FF",
	x"00", x"01", x"01", x"02", x"02", x"00", x"FF", x"FE", x"FE", x"FE", x"FD", x"FC",
	x"FB", x"FC", x"FC", x"FD", x"FE", x"00", x"02", x"02", x"02", x"02", x"03", x"03",
	x"02", x"01", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"00",
	x"01", x"02", x"01", x"FE", x"FD", x"FC", x"FD", x"FD", x"FC", x"FD", x"FE", x"FF",
	x"FF", x"00", x"01", x"01", x"03", x"02", x"01", x"01", x"00", x"00", x"00", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"02", x"01", x"00", x"FF",
	x"FF", x"FE", x"FD", x"FC", x"FD", x"FE", x"FE", x"FE", x"FF", x"00", x"02", x"02",
	x"01", x"02", x"01", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FE", x"FE", x"00",
	x"00", x"02", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FD", x"FD",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"01", x"02", x"01", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"00", x"02",
	x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FE", x"FE", x"FE", x"00",
	x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FE",
	x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FF",
	x"FE", x"FD", x"FF", x"FF", x"00", x"FF", x"FF", x"01", x"01", x"02", x"01", x"00",
	x"01", x"00", x"FF", x"FE", x"FF", x"FF", x"FE", x"FE", x"FD", x"FE", x"00", x"01",
	x"01", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"01", x"00", x"01", x"01", x"01", x"01", x"00", x"01", x"FE", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FE", x"FF", x"00", x"FF", x"01", x"03", x"03", x"02", x"01",
	x"00", x"FF", x"00", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"00",
	x"01", x"00", x"00", x"01", x"00", x"00", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"00", x"01", x"01", x"02", x"01", x"01", x"00", x"FF", x"FF",
	x"00", x"FF", x"FF", x"01", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF",
	x"FE", x"FD", x"FD", x"FE", x"FD", x"FC", x"FD", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"01", x"01", x"02", x"03", x"02", x"01", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FE", x"FD", x"FD", x"FD",
	x"FC", x"FD", x"FE", x"FF", x"00", x"00", x"02", x"03", x"03", x"02", x"02", x"02",
	x"02", x"01", x"00", x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"00", x"01", x"00", x"01", x"00", x"01", x"02", x"01",
	x"00", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"FE", x"FE", x"FD",
	x"FD", x"FD", x"FD", x"FB", x"FB", x"FD", x"FE", x"FF", x"00", x"02", x"03", x"03",
	x"02", x"03", x"03", x"02", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FD", x"FC", x"FD", x"FD", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"00", x"01", x"02", x"03", x"03", x"03", x"02", x"01", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"01",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FF", x"FF", x"00", x"01",
	x"01", x"02", x"03", x"02", x"01", x"01", x"01", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FD",
	x"FC", x"FC", x"FC", x"FC", x"FE", x"00", x"00", x"00", x"02", x"04", x"04", x"04",
	x"04", x"04", x"02", x"FF", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"00", x"02", x"02", x"02", x"03", x"01", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FD", x"FD", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"01", x"00", x"00", x"FF", x"FD", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"01",
	x"02", x"01", x"01", x"02", x"01", x"01", x"00", x"FE", x"FF", x"FF", x"FF", x"FD",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FE", x"FE", x"FD", x"FD",
	x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"02", x"01", x"02", x"02", x"01", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00",
	x"01", x"01", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"00", x"01", x"02", x"02", x"01", x"01", x"01", x"FF", x"FF", x"FF", x"FE", x"FD",
	x"FD", x"FE", x"FE", x"FF", x"01", x"00", x"00", x"00", x"01", x"01", x"00", x"FF",
	x"FF", x"FF", x"FD", x"FD", x"FF", x"00", x"00", x"01", x"00", x"00", x"00", x"01",
	x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF",
	x"00", x"00", x"00", x"01", x"02", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"02", x"01", x"00", x"FF", x"FF",
	x"FE", x"FC", x"FC", x"FC", x"FD", x"FE", x"FF", x"00", x"01", x"01", x"02", x"02",
	x"02", x"01", x"01", x"02", x"01", x"FF", x"FE", x"FE", x"FF", x"FE", x"FF", x"00",
	x"01", x"00", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"FE", x"FD", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"02", x"03", x"02", x"03", x"01",
	x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"FE", x"FC", x"FD", x"FD", x"FE", x"FE", x"FD", x"FE", x"FF", x"01", x"02",
	x"02", x"03", x"03", x"02", x"01", x"01", x"01", x"01", x"01", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FE", x"FD", x"FE", x"FF", x"00", x"01", x"02", x"02", x"02", x"02",
	x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE", x"00",
	x"00", x"FE", x"00", x"00", x"01", x"03", x"03", x"02", x"00", x"00", x"00", x"01",
	x"01", x"00", x"01", x"01", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FD",
	x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FD", x"FF", x"FF", x"00", x"02", x"04",
	x"05", x"04", x"04", x"04", x"02", x"03", x"01", x"FE", x"FD", x"FE", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FE", x"FD", x"FF", x"00", x"FF", x"FE", x"FD", x"FD",
	x"FD", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"02", x"03", x"03",
	x"02", x"01", x"00", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"01", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FC", x"FE", x"FE", x"FF",
	x"FF", x"01", x"02", x"03", x"04", x"04", x"03", x"02", x"02", x"00", x"00", x"00",
	x"FF", x"FE", x"FD", x"FD", x"FE", x"00", x"01", x"FF", x"FE", x"FE", x"FE", x"FD",
	x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FF", x"01", x"02", x"02", x"02", x"02",
	x"02", x"03", x"03", x"03", x"02", x"01", x"FE", x"FD", x"FC", x"FD", x"FD", x"FD",
	x"FE", x"FD", x"FE", x"00", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"00", x"01", x"02", x"02", x"02", x"01", x"00", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"02", x"00",
	x"01", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FE",
	x"00", x"03", x"03", x"02", x"01", x"02", x"01", x"01", x"00", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"00", x"FE",
	x"FD", x"FE", x"FD", x"FE", x"00", x"01", x"01", x"02", x"03", x"02", x"02", x"02",
	x"02", x"01", x"FF", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"01", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"02", x"01", x"01", x"00", x"01", x"00", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FD", x"FD", x"FF", x"00", x"01", x"02", x"01", x"01", x"02",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"00", x"01", x"02", x"02",
	x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FD", x"FC", x"FE",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"01", x"01", x"00", x"00",
	x"FF", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00",
	x"FF", x"FE", x"FD", x"FD", x"FE", x"FD", x"FD", x"FD", x"FD", x"FF", x"00", x"02",
	x"04", x"03", x"02", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FE", x"FE",
	x"FE", x"FE", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01",
	x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00",
	x"00", x"FF", x"00", x"00", x"FE", x"FD", x"FE", x"FD", x"FD", x"FE", x"FE", x"00",
	x"01", x"00", x"00", x"02", x"03", x"02", x"02", x"01", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FE", x"FD", x"FE", x"FF", x"FE", x"FD", x"FE", x"FF", x"FF", x"01", x"01", x"02",
	x"02", x"02", x"02", x"01", x"01", x"01", x"00", x"00", x"FE", x"FE", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FE", x"FD", x"FC",
	x"FD", x"FF", x"01", x"02", x"02", x"01", x"03", x"03", x"01", x"02", x"02", x"01",
	x"01", x"FF", x"FE", x"FE", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"00", x"00",
	x"01", x"03", x"03", x"04", x"04", x"03", x"02", x"02", x"00", x"FE", x"FE", x"FE",
	x"FD", x"FC", x"FD", x"FE", x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"01", x"02", x"02", x"02", x"02", x"01",
	x"01", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00",
	x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FD", x"FE", x"FD", x"FE", x"FF",
	x"FF", x"00", x"00", x"01", x"02", x"03", x"05", x"03", x"03", x"02", x"01", x"FF",
	x"FE", x"FE", x"FE", x"FD", x"FC", x"FC", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"01", x"01", x"01",
	x"01", x"02", x"02", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FD", x"FD",
	x"FD", x"FE", x"FE", x"FE", x"FF", x"01", x"01", x"00", x"FF", x"00", x"00", x"FF",
	x"FE", x"FD", x"FF", x"FF", x"00", x"01", x"00", x"01", x"02", x"02", x"00", x"01",
	x"01", x"01", x"00", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FE", x"FE", x"00", x"00",
	x"00", x"01", x"02", x"02", x"02", x"03", x"03", x"02", x"02", x"00", x"FF", x"FF",
	x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"02", x"02", x"03", x"03",
	x"02", x"01", x"00", x"FF", x"FF", x"FE", x"FD", x"FC", x"FC", x"FD", x"FD", x"FF",
	x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FD",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FE", x"FE", x"FE", x"FF", x"01", x"00", x"00",
	x"01", x"01", x"00", x"FE", x"FE", x"FD", x"FF", x"FF", x"FE", x"FF", x"FF", x"00",
	x"02", x"03", x"02", x"02", x"03", x"01", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD",
	x"FD", x"FD", x"FF", x"FF", x"00", x"00", x"01", x"02", x"01", x"01", x"00", x"00",
	x"01", x"00", x"FE", x"FE", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"01", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FD", x"FF", x"FF", x"FE", x"FF", x"00",
	x"01", x"01", x"02", x"02", x"02", x"01", x"01", x"00", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"00", x"01", x"01",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"01", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FD", x"FD", x"FD",
	x"FE", x"00", x"00", x"01", x"01", x"02", x"02", x"01", x"02", x"02", x"01", x"00",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FF", x"00", x"FE", x"FE", x"FF", x"00", x"FF", x"00", x"01", x"00", x"01", x"02",
	x"01", x"01", x"02", x"02", x"02", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FD",
	x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FE", x"FD", x"FE", x"FF",
	x"FE", x"FE", x"FE", x"FF", x"01", x"02", x"01", x"03", x"05", x"03", x"02", x"02",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE", x"FE", x"FD", x"FE", x"FF", x"00",
	x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"00", x"01", x"02", x"02", x"03", x"04", x"03", x"03", x"02", x"00", x"FF", x"FF",
	x"FE", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"01", x"00", x"01", x"02", x"02", x"02",
	x"03", x"02", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FF", x"FF", x"00", x"00", x"01", x"03", x"04", x"03", x"02", x"01", x"01",
	x"01", x"00", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FD", x"FE", x"00", x"00", x"01",
	x"01", x"02", x"01", x"01", x"01", x"01", x"01", x"01", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FF",
	x"FE", x"FE", x"FF", x"FD", x"FE", x"FE", x"00", x"01", x"01", x"03", x"03", x"02",
	x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FD", x"FD", x"FF", x"FF",
	x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"01", x"02", x"02", x"02", x"02", x"02", x"01", x"01", x"00", x"FE",
	x"FF", x"FF", x"FE", x"FC", x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"FF",
	x"01", x"02", x"01", x"02", x"01", x"00", x"FF", x"FE", x"FD", x"FE", x"FF", x"FE",
	x"FE", x"00", x"00", x"00", x"02", x"02", x"02", x"01", x"00", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01",
	x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"00", x"00",
	x"00", x"02", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FD",
	x"FD", x"FE", x"FE", x"FF", x"01", x"01", x"01", x"01", x"01", x"01", x"02", x"02",
	x"01", x"00", x"FF", x"FE", x"FD", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FF",
	x"FF", x"FF", x"00", x"01", x"00", x"00", x"FF", x"FF", x"00", x"01", x"00", x"FF",
	x"01", x"02", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FD", x"FD", x"FD", x"FD", x"FF", x"01", x"00", x"00", x"01", x"01", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"01", x"01", x"01", x"00", x"01",
	x"01", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FD", x"FD", x"FD",
	x"FE", x"FE", x"FE", x"00", x"01", x"01", x"02", x"03", x"04", x"03", x"02", x"01",
	x"00", x"FF", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01",
	x"01", x"02", x"03", x"02", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FD",
	x"FD", x"FD", x"FE", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"02", x"02", x"02",
	x"03", x"02", x"01", x"00", x"FE", x"FD", x"FD", x"FE", x"FD", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"00",
	x"00", x"00", x"01", x"01", x"01", x"01", x"02", x"03", x"03", x"02", x"00", x"FF",
	x"00", x"FF", x"FD", x"FD", x"FC", x"FC", x"FD", x"FE", x"FE", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"01", x"01", x"00", x"FE", x"FF", x"00", x"01", x"02", x"02",
	x"02", x"01", x"01", x"00", x"FF", x"FF", x"00", x"FF", x"FD", x"FC", x"FD", x"FE",
	x"FF", x"FF", x"00", x"01", x"01", x"FF", x"00", x"01", x"00", x"FF", x"00", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"02", x"02",
	x"01", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF",
	x"00", x"01", x"00", x"00", x"FF", x"FE", x"FF", x"00", x"FF", x"FE", x"FF", x"00",
	x"FF", x"00", x"02", x"02", x"03", x"03", x"02", x"FF", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FD", x"FF", x"01", x"01", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"01", x"02", x"02",
	x"01", x"01", x"02", x"01", x"00", x"FF", x"FD", x"FC", x"FD", x"FE", x"FE", x"FE",
	x"00", x"FF", x"00", x"01", x"01", x"02", x"02", x"01", x"FF", x"FE", x"FD", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"02", x"02", x"02", x"01", x"FF",
	x"FE", x"FD", x"FE", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"01",
	x"02", x"01", x"01", x"00", x"FF", x"00", x"FF", x"FD", x"FD", x"FE", x"FF", x"FF",
	x"FF", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FD",
	x"FD", x"FE", x"FF", x"00", x"00", x"02", x"02", x"01", x"01", x"01", x"01", x"00",
	x"FF", x"FE", x"FD", x"FD", x"FD", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"01", x"02", x"01", x"00", x"FF", x"FE", x"FF", x"FF", x"FD", x"FD",
	x"FE", x"FE", x"FE", x"FE", x"00", x"01", x"02", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"03", x"03", x"01", x"01",
	x"01", x"00", x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"01", x"00", x"00", x"01", x"01", x"00",
	x"00", x"00", x"01", x"01", x"01", x"00", x"FF", x"00", x"00", x"FF", x"FE", x"FD",
	x"FD", x"FD", x"FE", x"FF", x"FE", x"FE", x"00", x"00", x"FF", x"00", x"01", x"02",
	x"01", x"FF", x"FE", x"FD", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"02", x"01",
	x"02", x"03", x"03", x"01", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FD", x"FE",
	x"FD", x"FD", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"01", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"01", x"02", x"02", x"02", x"02", x"02", x"02", x"02",
	x"01", x"01", x"FF", x"FC", x"FC", x"FC", x"FC", x"FC", x"FD", x"FD", x"FD", x"FE",
	x"FF", x"FF", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"02",
	x"02", x"03", x"01", x"01", x"02", x"01", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD",
	x"FC", x"FC", x"FE", x"FD", x"FE", x"FE", x"FF", x"01", x"01", x"01", x"00", x"01",
	x"01", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"01", x"03", x"03",
	x"03", x"02", x"01", x"00", x"01", x"00", x"FE", x"FD", x"FC", x"FB", x"FB", x"FC",
	x"FD", x"FE", x"00", x"FF", x"FE", x"FF", x"00", x"01", x"01", x"00", x"00", x"01",
	x"01", x"00", x"01", x"02", x"02", x"02", x"01", x"01", x"00", x"00", x"01", x"FF",
	x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FC", x"FD", x"FE", x"FE", x"FF", x"00",
	x"01", x"01", x"01", x"00", x"FF", x"00", x"01", x"01", x"00", x"00", x"00", x"00",
	x"01", x"00", x"01", x"02", x"01", x"00", x"FF", x"FE", x"FE", x"FD", x"FE", x"FD",
	x"FD", x"FE", x"FE", x"FF", x"FF", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"01", x"02", x"02", x"01",
	x"02", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"00", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF",
	x"01", x"02", x"02", x"02", x"01", x"01", x"03", x"02", x"01", x"00", x"FF", x"FE",
	x"FC", x"FB", x"FC", x"FD", x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"02", x"02",
	x"01", x"01", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"00", x"01",
	x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FD",
	x"FD", x"FF", x"00", x"01", x"01", x"01", x"01", x"02", x"01", x"01", x"00", x"FF",
	x"FE", x"FD", x"FD", x"FD", x"FE", x"FF", x"00", x"01", x"01", x"02", x"01", x"01",
	x"01", x"00", x"00", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF", x"00", x"01", x"00",
	x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"02", x"02", x"02", x"02", x"00",
	x"00", x"00", x"FE", x"FE", x"FE", x"FC", x"FC", x"FD", x"FE", x"FE", x"00", x"01",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01",
	x"02", x"02", x"01", x"01", x"01", x"01", x"00", x"00", x"FE", x"FE", x"FE", x"FD",
	x"FC", x"FD", x"FE", x"FE", x"FF", x"FE", x"FF", x"01", x"01", x"01", x"01", x"01",
	x"00", x"FF", x"FF", x"FE", x"FE", x"00", x"01", x"00", x"01", x"02", x"01", x"02",
	x"02", x"02", x"01", x"00", x"FF", x"FD", x"FC", x"FD", x"FD", x"FE", x"FF", x"FE",
	x"FE", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"01",
	x"00", x"00", x"02", x"01", x"02", x"03", x"02", x"01", x"01", x"01", x"FF", x"FF",
	x"FF", x"FE", x"FD", x"FC", x"FC", x"FD", x"FD", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"00", x"00", x"01", x"02",
	x"03", x"03", x"03", x"03", x"03", x"02", x"00", x"FF", x"FE", x"FD", x"FC", x"FB",
	x"FC", x"FC", x"FC", x"FD", x"FE", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"02", x"02", x"02", x"02",
	x"01", x"00", x"FF", x"FF", x"FE", x"FD", x"FD", x"FC", x"FC", x"FB", x"FC", x"FD",
	x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"02", x"03", x"02", x"02", x"02", x"01", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FD", x"FC", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01",
	x"02", x"02", x"02", x"02", x"01", x"01", x"00", x"FE", x"FD", x"FE", x"FD", x"FC",
	x"FC", x"FC", x"FC", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"00",
	x"01", x"01", x"01", x"01", x"02", x"02", x"01", x"01", x"01", x"01", x"00", x"FF",
	x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FF", x"FF", x"00",
	x"01", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF",
	x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"02", x"01", x"00", x"FE", x"FD",
	x"FC", x"FC", x"FD", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"00",
	x"00", x"FF", x"FD", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"01", x"03", x"02",
	x"02", x"02", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FD", x"FC", x"FC", x"FC",
	x"FD", x"FF", x"00", x"00", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"00",
	x"FF", x"FF", x"FF", x"00", x"01", x"00", x"01", x"01", x"01", x"00", x"00", x"FF",
	x"FE", x"FE", x"FD", x"FC", x"FC", x"FD", x"FD", x"FF", x"00", x"01", x"02", x"03",
	x"02", x"02", x"02", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"00", x"00", x"00", x"01", x"02", x"01", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"00",
	x"00", x"01", x"02", x"01", x"01", x"02", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FE", x"FE", x"00", x"00", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"02", x"02", x"01", x"01", x"01",
	x"01", x"00", x"00", x"FF", x"FD", x"FD", x"FD", x"FC", x"FE", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FF", x"00", x"00",
	x"00", x"01", x"01", x"01", x"01", x"02", x"01", x"00", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FD", x"FD", x"FF", x"00", x"FF", x"00", x"01", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01",
	x"02", x"02", x"02", x"02", x"02", x"01", x"00", x"FE", x"FE", x"FD", x"FC", x"FD",
	x"FE", x"FE", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"00", x"00", x"00", x"01", x"02", x"02", x"03", x"03", x"02", x"02", x"02", x"00",
	x"FF", x"FE", x"FE", x"FD", x"FD", x"FC", x"FC", x"FD", x"FE", x"FE", x"FE", x"FF",
	x"01", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"00", x"01", x"03", x"03", x"03", x"02", x"00", x"FF", x"FF", x"FE", x"FD",
	x"FC", x"FD", x"FD", x"FC", x"FD", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00",
	x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FD",
	x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"01", x"01", x"FF", x"FF", x"00",
	x"00", x"01", x"01", x"02", x"02", x"02", x"01", x"01", x"01", x"01", x"00", x"FF",
	x"FD", x"FD", x"FC", x"FC", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"01",
	x"01", x"01", x"01", x"01", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FD",
	x"FC", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"02",
	x"00", x"00", x"00", x"FF", x"FF", x"01", x"02", x"02", x"02", x"01", x"01", x"01",
	x"00", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FD", x"FF", x"FF", x"FE",
	x"FF", x"01", x"01", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"01", x"02", x"02", x"01", x"01", x"01", x"00", x"FF",
	x"FF", x"FD", x"FD", x"FD", x"FC", x"FC", x"FD", x"FE", x"FF", x"00", x"01", x"00",
	x"01", x"01", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"02",
	x"02", x"02", x"02", x"00", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FC", x"FD",
	x"FD", x"FD", x"FE", x"00", x"01", x"00", x"01", x"02", x"02", x"02", x"01", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"02",
	x"01", x"FF", x"FE", x"FE", x"FD", x"FE", x"FF", x"FE", x"FE", x"FF", x"00", x"00",
	x"01", x"02", x"02", x"02", x"01", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FE", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"FF", x"00", x"01", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"00", x"00",
	x"00", x"01", x"01", x"00", x"FF", x"00", x"FF", x"FD", x"FC", x"FD", x"FE", x"FF",
	x"00", x"01", x"01", x"02", x"02", x"02", x"02", x"01", x"FF", x"FF", x"FE", x"FD",
	x"FD", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"FF", x"00", x"01", x"02", x"01",
	x"01", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"FF",
	x"00", x"01", x"01", x"02", x"02", x"01", x"00", x"00", x"01", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"02", x"01", x"01", x"01", x"00", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"01", x"01",
	x"01", x"01", x"02", x"01", x"02", x"02", x"00", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FD", x"FD", x"FC", x"FC", x"FE", x"FF", x"01", x"01", x"01", x"01", x"00", x"FF",
	x"FF", x"00", x"01", x"00", x"01", x"00", x"01", x"03", x"02", x"01", x"01", x"00",
	x"FF", x"FF", x"FE", x"FD", x"FE", x"FE", x"FC", x"FB", x"FC", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"01", x"01", x"02", x"02", x"02", x"01", x"00", x"00", x"FE", x"FF",
	x"00", x"01", x"00", x"FF", x"00", x"00", x"00", x"01", x"02", x"01", x"00", x"00",
	x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FD", x"FD", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"02", x"02", x"01", x"01", x"01",
	x"01", x"00", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FD", x"FC", x"FD",
	x"FD", x"FD", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"02", x"01",
	x"01", x"00", x"FF", x"FF", x"00", x"00", x"01", x"02", x"01", x"00", x"00", x"01",
	x"00", x"00", x"FF", x"FD", x"FC", x"FC", x"FD", x"FD", x"FE", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"00", x"01", x"01", x"FF",
	x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"00", x"FF", x"FF", x"01", x"01", x"00", x"FF", x"00", x"00", x"01", x"02", x"01",
	x"02", x"02", x"01", x"FF", x"FF", x"FE", x"FD", x"FE", x"FD", x"FC", x"FC", x"FE",
	x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"01", x"00", x"FF",
	x"FF", x"FE", x"FF", x"01", x"01", x"FF", x"00", x"01", x"01", x"01", x"01", x"01",
	x"00", x"FF", x"FE", x"FC", x"FD", x"FE", x"FE", x"FE", x"FD", x"FD", x"FF", x"00",
	x"01", x"01", x"02", x"02", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"01", x"01",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"00", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"00", x"00", x"00", x"FF", x"00", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FD",
	x"FD", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"02", x"01", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"01", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FE", x"FD", x"FE", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FE", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"FF", x"FF", x"FF",
	x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"02", x"01",
	x"01", x"00", x"01", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FE", x"FF",
	x"FF", x"FF", x"00", x"00", x"01", x"03", x"03", x"02", x"01", x"00", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"00", x"01", x"01", x"02", x"02", x"01",
	x"00", x"00", x"FF", x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"FF", x"00", x"00", x"00", x"01",
	x"02", x"02", x"01", x"01", x"00", x"FF", x"01", x"01", x"FF", x"FE", x"FD", x"FC",
	x"FC", x"FC", x"FD", x"FD", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"02", x"02",
	x"02", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"01", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FE", x"FD", x"FD", x"FE", x"FD", x"FE", x"FF", x"FF",
	x"FF", x"00", x"01", x"00", x"01", x"01", x"00", x"00", x"00", x"01", x"01", x"01",
	x"00", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"00", x"FF",
	x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"01", x"01", x"01",
	x"02", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FC", x"FC", x"FD", x"FD",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"02", x"02", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FD", x"FE", x"FF", x"00", x"00", x"00",
	x"01", x"00", x"FF", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FF", x"00",
	x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"00", x"01", x"00", x"00", x"FF",
	x"FF", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"01",
	x"01", x"02", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FE", x"FF", x"00", x"02", x"02", x"02", x"02", x"01", x"01", x"00", x"00",
	x"FF", x"FF", x"FE", x"FD", x"FE", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"01", x"00", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF",
	x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"02", x"01", x"01", x"01",
	x"00", x"FF", x"FE", x"FF", x"FF", x"FE", x"FF", x"FE", x"FE", x"FE", x"FF", x"00",
	x"01", x"01", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FE", x"FF", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FF",
	x"FE", x"FD", x"FD", x"FE", x"FF", x"00", x"01", x"01", x"01", x"02", x"02", x"01",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"01", x"00", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FD", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"00", x"FF",
	x"FE", x"FD", x"FD", x"FE", x"FD", x"FD", x"FE", x"FF", x"00", x"01", x"02", x"01",
	x"02", x"02", x"00", x"00", x"01", x"00", x"FE", x"FF", x"FE", x"FE", x"FF", x"00",
	x"00", x"01", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FD", x"FD",
	x"FE", x"FE", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"02", x"02", x"01",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"01", x"02",
	x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FD", x"FC", x"FC", x"FD", x"FE", x"FF",
	x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"00", x"00", x"00", x"01", x"00", x"FF", x"FE", x"FE", x"FD", x"FD", x"FD",
	x"FD", x"FE", x"FD", x"FD", x"FD", x"FE", x"00", x"00", x"01", x"03", x"03", x"03",
	x"02", x"02", x"02", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"FF",
	x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00",
	x"FF", x"FE", x"FD", x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"FF", x"00", x"00",
	x"01", x"01", x"01", x"02", x"02", x"02", x"01", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FD", x"FC", x"FD",
	x"FD", x"FD", x"FE", x"FF", x"00", x"01", x"02", x"02", x"02", x"02", x"02", x"02",
	x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"00", x"01", x"01", x"00", x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"00", x"01", x"00", x"FF", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"01", x"02", x"00", x"00", x"00", x"FF", x"FE",
	x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"00", x"00", x"00", x"01",
	x"02", x"02", x"02", x"02", x"02", x"02", x"01", x"FF", x"FF", x"FF", x"FD", x"FE",
	x"FF", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FE",
	x"FE", x"FF", x"FE", x"FE", x"00", x"01", x"01", x"02", x"02", x"01", x"01", x"02",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"00",
	x"01", x"00", x"00", x"01", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FE",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"00",
	x"FF", x"FE", x"FE", x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"01",
	x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FF", x"00", x"00", x"00", x"01", x"02", x"03",
	x"03", x"02", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00",
	x"00", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FD", x"FD", x"FE",
	x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"01", x"01", x"00",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FD", x"FD", x"FD", x"FC", x"FD", x"FE", x"FF", x"00", x"02",
	x"01", x"02", x"02", x"01", x"01", x"01", x"01", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FD",
	x"FD", x"FD", x"FE", x"FD", x"FE", x"FF", x"FF", x"01", x"02", x"02", x"02", x"02",
	x"01", x"00", x"01", x"00", x"00", x"01", x"00", x"FE", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE",
	x"FF", x"00", x"00", x"01", x"02", x"02", x"01", x"01", x"02", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FE", x"FE",
	x"FD", x"FC", x"FC", x"FD", x"FD", x"FE", x"FF", x"00", x"00", x"01", x"01", x"02",
	x"03", x"03", x"03", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE",
	x"FD", x"FE", x"00", x"00", x"FF", x"00", x"01", x"02", x"01", x"01", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FD", x"FD", x"FE", x"FF", x"00", x"01",
	x"01", x"01", x"02", x"02", x"02", x"02", x"02", x"02", x"00", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FE",
	x"FE", x"FD", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"03", x"03", x"01",
	x"02", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"02", x"01", x"01", x"01", x"01",
	x"01", x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"00", x"01", x"01", x"01",
	x"02", x"02", x"03", x"03", x"03", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FD", x"FE", x"FD", x"FC", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01",
	x"02", x"02", x"01", x"01", x"00", x"FE", x"FD", x"FD", x"FE", x"FD", x"FD", x"FD",
	x"FE", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"01", x"00",
	x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE", x"FF", x"00", x"00", x"01", x"02",
	x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FD", x"FD", x"FE", x"FF",
	x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"FF", x"00", x"01", x"01", x"01",
	x"01", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FD", x"FE",
	x"00", x"01", x"02", x"03", x"02", x"02", x"02", x"01", x"01", x"00", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FE",
	x"FE", x"FD", x"FD", x"FD", x"FE", x"FF", x"00", x"00", x"00", x"00", x"01", x"02",
	x"02", x"02", x"01", x"01", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"00", x"01", x"01", x"02", x"02", x"02", x"02", x"01", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"00", x"00", x"FE",
	x"FD", x"FD", x"FD", x"FD", x"FE", x"FE", x"FD", x"FE", x"FF", x"00", x"02", x"02",
	x"02", x"02", x"02", x"01", x"01", x"01", x"02", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"01", x"02", x"02", x"01",
	x"01", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FD", x"FC", x"FD", x"FE", x"FE", x"FF", x"FF",
	x"00", x"00", x"01", x"02", x"03", x"02", x"01", x"01", x"01", x"01", x"00", x"00",
	x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"01", x"02", x"02", x"02", x"01", x"00", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"FF", x"FE", x"FD", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"02", x"02", x"02", x"02",
	x"01", x"00", x"01", x"00", x"FF", x"FF", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FD", x"FE", x"FF", x"00", x"01",
	x"02", x"03", x"02", x"02", x"01", x"02", x"01", x"00", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FE", x"FF", x"00", x"01", x"02", x"02", x"02", x"01", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"01", x"01", x"00", x"01", x"01", x"00", x"FE", x"FD", x"FD", x"FE", x"FE",
	x"FE", x"FF", x"00", x"01", x"01", x"01", x"02", x"02", x"02", x"01", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01",
	x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"01", x"02", x"01", x"01", x"01", x"01", x"01", x"FF", x"FE",
	x"FE", x"FE", x"FC", x"FD", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"FF", x"FF", x"00", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FE", x"FD", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"02", x"03", x"03", x"03", x"02", x"01", x"01", x"00",
	x"FE", x"FD", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01",
	x"01", x"01", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"01", x"00", x"FE", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"02", x"02", x"02", x"01",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"01", x"01", x"02", x"03", x"02", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01",
	x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FF", x"00", x"00", x"00", x"01", x"01", x"02", x"02", x"02", x"02", x"02", x"01",
	x"00", x"FF", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"00",
	x"01", x"02", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"00", x"01", x"01", x"00", x"00",
	x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"01", x"02", x"01", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"00", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"02", x"02", x"02", x"01", x"00",
	x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FE", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"01", x"02", x"02", x"02",
	x"02", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"01", x"02", x"02", x"02", x"02", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FD", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"01", x"01", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"01",
	x"00", x"00", x"01", x"01", x"00", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"02", x"02", x"02", x"02",
	x"01", x"01", x"00", x"FF", x"FE", x"FD", x"FD", x"FE", x"FD", x"FD", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"01", x"02", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"01", x"01", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"02", x"02", x"02", x"02", x"01", x"01",
	x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"01", x"00", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"01", x"00", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"01",
	x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"02", x"01",
	x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FF",
	x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"FF", x"00", x"01", x"01", x"01", x"00", x"01", x"00", x"00", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"02", x"02",
	x"02", x"02", x"02", x"02", x"01", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"01", x"01", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"00", x"01", x"01", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00",
	x"01", x"02", x"02", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FD",
	x"FD", x"FD", x"FE", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"00", x"01", x"02", x"02", x"02", x"02", x"02",
	x"02", x"01", x"01", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FC", x"FD", x"FD",
	x"FD", x"FE", x"00", x"00", x"01", x"00", x"00", x"01", x"01", x"00", x"00", x"01",
	x"00", x"FF", x"00", x"00", x"00", x"01", x"02", x"01", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"01", x"02", x"01", x"00", x"00", x"01", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"01", x"02", x"02",
	x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FE", x"FD", x"FD", x"FD", x"FE",
	x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"01", x"00",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FD", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"01", x"01",
	x"02", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"01", x"01", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"00", x"00",
	x"01", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"00", x"00", x"01", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01",
	x"02", x"02", x"01", x"01", x"01", x"FF", x"FE", x"FD", x"FD", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"02", x"02", x"02", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FC", x"FC",
	x"FC", x"FC", x"FD", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"01", x"02", x"02", x"01", x"00", x"01",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"02", x"03", x"02", x"02", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FD", x"FD", x"FD", x"FC", x"FD", x"FF", x"00", x"00", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"02", x"02",
	x"02", x"02", x"02", x"01", x"00", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD",
	x"FD", x"FD", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"FF",
	x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00",
	x"FF", x"FF", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"01", x"02", x"02", x"02", x"02", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FE",
	x"FD", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"FF", x"00", x"02", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00",
	x"01", x"02", x"02", x"02", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FD",
	x"FD", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"01", x"02", x"02", x"02", x"01", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"01", x"01", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"01", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FD", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"02", x"01", x"01", x"00", x"00",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"01", x"01", x"01",
	x"02", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FD", x"FD", x"FD",
	x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"01", x"02", x"02", x"01", x"01", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"00", x"01",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"01", x"01", x"01", x"02", x"02", x"02", x"01", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FD", x"FE", x"FD", x"FC", x"FD", x"FE", x"FF", x"01", x"02", x"01", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"02", x"02", x"02",
	x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE",
	x"FE", x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"01", x"01", x"00", x"01", x"01", x"02", x"01", x"01", x"01", x"00",
	x"FF", x"FD", x"FC", x"FC", x"FD", x"FE", x"FD", x"FE", x"FF", x"00", x"00", x"00",
	x"00", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01",
	x"01", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FD", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"01",
	x"01", x"01", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"01", x"02", x"02", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FD", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF", x"00",
	x"00", x"00", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"01", x"02", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"00", x"00", x"00", x"01", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01",
	x"00", x"00", x"00", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"02", x"02", x"01", x"00", x"00",
	x"00", x"00", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"01", x"00", x"00", x"00", x"01", x"00", x"00", x"01",
	x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FD",
	x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01",
	x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"00", x"01", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"02", x"02", x"01", x"FF", x"FF",
	x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"01",
	x"02", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FD", x"FD", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"01", x"01", x"02", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FE", x"FD", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"FF", x"FF", x"FE", x"FF", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FE", x"FE", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"01", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"01", x"01", x"00",
	x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"01",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01",
	x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"01", x"01", x"02", x"01", x"01", x"01", x"00", x"FF", x"00", x"01", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FE", x"FF",
	x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FF", x"FE", x"FD", x"FE", x"FE", x"FF", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FF", x"00",
	x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01",
	x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FD",
	x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"02", x"01", x"01",
	x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FD", x"FE", x"FF",
	x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"FE",
	x"FD", x"FD", x"FD", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"00", x"01", x"01",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"01", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"00",
	x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"01", x"02", x"02", x"01", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"01", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FE", x"FF", x"00",
	x"01", x"01", x"01", x"02", x"02", x"02", x"02", x"01", x"00", x"00", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"02", x"02", x"02",
	x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD",
	x"FD", x"FE", x"FF", x"00", x"01", x"02", x"01", x"01", x"01", x"02", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FD", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"01", x"02", x"01", x"01", x"01", x"00", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"00", x"FF", x"FE", x"FE", x"FD",
	x"FD", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"01", x"02", x"01", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE",
	x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"02", x"02", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"02", x"02", x"02",
	x"02", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"01", x"02", x"01",
	x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF", x"00", x"00",
	x"01", x"01", x"01", x"01", x"02", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01",
	x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"01", x"01", x"01", x"02", x"01", x"01", x"01", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"02", x"02", x"01", x"01", x"00", x"FF", x"FF", x"00", x"FF", x"FE", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"02", x"02", x"02", x"02",
	x"01", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"01", x"01", x"01", x"01", x"01", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"00", x"01", x"02", x"02", x"02",
	x"02", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"00", x"01", x"01", x"02", x"01", x"01", x"01", x"01", x"00", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"02",
	x"02", x"02", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01",
	x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FD", x"FD", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00",
	x"00", x"01", x"02", x"02", x"02", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01",
	x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF",
	x"FF", x"FE", x"FF", x"00", x"00", x"00", x"01", x"01", x"02", x"02", x"02", x"01",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00",
	x"01", x"01", x"02", x"02", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"01", x"01",
	x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"FF",
	x"00", x"00", x"01", x"02", x"03", x"02", x"01", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"00", x"01", x"02",
	x"02", x"02", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"01", x"01", x"01",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00",
	x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"02", x"02", x"01", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"02", x"02", x"02", x"01",
	x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"02", x"02", x"01", x"01", x"00", x"01",
	x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FD", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FD", x"FE", x"FE", x"FD", x"FE", x"FE",
	x"FF", x"00", x"01", x"02", x"02", x"02", x"02", x"02", x"01", x"01", x"00", x"00",
	x"FF", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"01", x"01", x"01", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"01", x"01", x"01", x"00", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"01",
	x"01", x"02", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"01", x"01", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE",
	x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"01", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"01", x"02", x"02", x"02", x"02", x"01", x"01", x"00",
	x"FF", x"FF", x"FE", x"FD", x"FD", x"FC", x"FD", x"FD", x"FF", x"00", x"00", x"01",
	x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"01", x"02",
	x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01",
	x"01", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FF", x"FF", x"00",
	x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01",
	x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"01",
	x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"02", x"01", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"01", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"01", x"02", x"02", x"02", x"01", x"01",
	x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01",
	x"02", x"02", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD",
	x"FD", x"FD", x"FD", x"FE", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"00", x"01", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"01",
	x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"00",
	x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"00", x"01", x"01", x"02", x"02", x"02", x"01", x"01", x"00", x"00", x"FF", x"FE",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00",
	x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"01", x"01",
	x"02", x"02", x"02", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FD",
	x"FD", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"01",
	x"01", x"00", x"00", x"00", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"01", x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FD", x"FD",
	x"FD", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01",
	x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01",
	x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FE", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"01", x"02", x"02", x"01", x"01", x"00", x"00", x"FF",
	x"FE", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"01", x"00", x"00", x"00", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"02", x"02", x"02", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"01", x"01", x"01", x"00", x"01", x"01", x"00", x"FE", x"FD", x"FD", x"FD",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00",
	x"FF", x"FE", x"FD", x"FD", x"FD", x"FE", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"00", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"02", x"01", x"01", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"00",
	x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"01", x"00",
	x"00", x"FF", x"FE", x"FE", x"FD", x"FE", x"FF", x"00", x"00", x"01", x"00", x"00",
	x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"01", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01",
	x"01", x"00", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"01", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FE", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"01",
	x"00", x"FF", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"00", x"01", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"01",
	x"01", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00",
	x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"01",
	x"01", x"01", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"01",
	x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"01",
	x"01", x"02", x"02", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"00", x"00", x"00", x"01", x"00", x"01", x"01", x"01", x"01", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01", x"00",
	x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"00",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF",
	x"00", x"01", x"01", x"01", x"02", x"02", x"02", x"02", x"01", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01",
	x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"01",
	x"00", x"00", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF",
	x"FF", x"FE", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"00", x"01", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01",
	x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"02", x"02", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"00", x"00", x"FF", x"00", x"01", x"01", x"01", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FD", x"FD", x"FE", x"00", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FE", x"FE", x"FD", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"01",
	x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"01", x"01", x"02", x"02",
	x"02", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FE", x"FE", x"FF",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00",
	x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"01", x"00", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"01", x"02", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FE",
	x"FE", x"FF", x"00", x"00", x"00", x"01", x"01", x"02", x"02", x"02", x"01", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FE", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"01", x"01", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"02", x"02", x"02",
	x"01", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FF", x"00", x"00", x"00",
	x"00", x"01", x"02", x"02", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"00", x"01", x"01", x"01", x"00", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"00", x"00", x"01", x"02", x"02", x"02", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01",
	x"00", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01",
	x"01", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FE", x"FE", x"FF",
	x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"01", x"01",
	x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FE",
	x"FE", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01",
	x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01",
	x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01",
	x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"00", x"01", x"01", x"01", x"02", x"01", x"01", x"01", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01",
	x"00", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"01",
	x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"FF", x"00",
	x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"01", x"00", x"00",
	x"01", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"01", x"02",
	x"02", x"02", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"01", x"01", x"02", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01",
	x"02", x"02", x"02", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FD", x"FD", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"01", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"02", x"02", x"01",
	x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FD", x"FD", x"FD", x"FE", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"01", x"02", x"02", x"02", x"02", x"01", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FE",
	x"FE", x"FD", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01",
	x"02", x"02", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"02", x"01", x"01", x"00", x"00",
	x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01",
	x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"01", x"02", x"02", x"01", x"01", x"01", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"02", x"01", x"01", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"01", x"02", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"02", x"02", x"01", x"01", x"00",
	x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01",
	x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"01", x"01", x"02", x"02", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01",
	x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01",
	x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"02", x"02", x"01",
	x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01",
	x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01",
	x"01", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF",
	x"FE", x"FE", x"FD", x"FD", x"FD", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"01",
	x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01",
	x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01",
	x"01", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FD", x"FD", x"FE", x"FF", x"00", x"01", x"01", x"01", x"01",
	x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FE", x"FE", x"FD", x"FD", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"01", x"02", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01",
	x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FD", x"FD", x"FE", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"01",
	x"02", x"02", x"02", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"00",
	x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"00",
	x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FE", x"FE", x"FE", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FD", x"FD", x"FD", x"FD", x"FE",
	x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01", x"02", x"02", x"01", x"01", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"01",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"01",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01",
	x"01", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"01", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00",
	x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"01", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01",
	x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01",
	x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00",
	x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01",
	x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"01", x"01", x"00", x"00",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01",
	x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01",
	x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"01", x"02", x"02", x"02", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"01", x"01", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00",
	x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"01",
	x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01",
	x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"01", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01",
	x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01",
	x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"01", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"00",
	x"00", x"00", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"01",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FE", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"01", x"01", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01",
	x"01", x"01", x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01",
	x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FE",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"00",
	x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01",
	x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01",
	x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01", x"01",
	x"01", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE",
	x"FE", x"FF", x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FE",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"01",
	x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FE", x"FE", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FE", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FE", x"FE", x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"01",
	x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FE",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00",
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"00", x"FF",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00",
	x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	x"FF", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"FF", x"FF",
	x"FF", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"FF", x"00",
	x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"00",
	x"00", x"FF", x"00", x"FF", x"FF", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF",
	x"00", x"FF", x"00", x"FF", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00",
	x"FF", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00",
	x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF",
	x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"00", x"00", x"00", x"00",
	x"00", x"00", x"00", x"FF", x"00", x"FF", x"00", x"FF", x"00", x"00", x"00", x"FF",
	x"FF", x"00", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00"
	);
	
signal cnt_out: unsigned(17 downto 0) := (others => '0');	
signal play_sound: std_logic := '0';
constant cnt_max: integer := 107519;
signal out_signal: signed(7 downto 0) := x"00";

begin
	
process (CLK)
begin
    if rising_edge(CLK) then
        if RST = '1' then
            play_sound <= '0';
        elsif PLAY = '1' then
            play_sound <= '1';
        elsif PLAY = '0' and cnt_out = cnt_max then
            play_sound <= '0';
        end if;
    end if;
end process;

	
-- 12bit counter
process (CLK)
begin     
    if rising_edge(CLK) then
        if RST = '1' then
            cnt_out <= (others => '0');
        elsif CE = '1' and play_sound = '1' then
            cnt_out <= cnt_out + 1;       
        end if;
        if cnt_out = cnt_max then
            cnt_out <= (others => '0');            
        end if;        
    end if;
end process;

--SAMPLE_OUT <= kick_sound(conv_integer(cnt_out));
process (CLK) 
begin
    if rising_edge(CLK) then
        if RST = '1' then
            out_signal <= x"00";
        elsif CE = '1' then
            out_signal <= ride_sound(conv_integer(cnt_out));
        end if;
    end if;    
end process;

SAMPLE_OUT <= out_signal;

end Behavioral;
